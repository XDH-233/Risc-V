// Generator : SpinalHDL v1.4.0    git head : ecb5a80b713566f417ea3ea061f9969e73770a7f
// Date      : 13/08/2021, 20:23:05
// Component : dataMem



module dataMem (
  input      [12:0]   address,
  input      [63:0]   writeData,
  output reg [63:0]   readData,
  input               memRead,
  input               memWrite,
  input               clk,
  input               reset 
);
  wire       [63:0]   _zz_2_;
  wire       [9:0]    _zz_3_;
  wire       [63:0]   content_0;
  wire       [63:0]   content_1;
  wire       [63:0]   content_2;
  wire       [63:0]   content_3;
  wire       [63:0]   content_4;
  wire       [63:0]   content_5;
  wire       [63:0]   content_6;
  wire       [63:0]   content_7;
  wire       [63:0]   content_8;
  wire       [63:0]   content_9;
  wire       [63:0]   content_10;
  wire       [63:0]   content_11;
  wire       [63:0]   content_12;
  wire       [63:0]   content_13;
  wire       [63:0]   content_14;
  wire       [63:0]   content_15;
  wire       [63:0]   content_16;
  wire       [63:0]   content_17;
  wire       [63:0]   content_18;
  wire       [63:0]   content_19;
  wire       [63:0]   content_20;
  wire       [63:0]   content_21;
  wire       [63:0]   content_22;
  wire       [63:0]   content_23;
  wire       [63:0]   content_24;
  wire       [63:0]   content_25;
  wire       [63:0]   content_26;
  wire       [63:0]   content_27;
  wire       [63:0]   content_28;
  wire       [63:0]   content_29;
  wire       [63:0]   content_30;
  wire       [63:0]   content_31;
  wire       [63:0]   content_32;
  wire       [63:0]   content_33;
  wire       [63:0]   content_34;
  wire       [63:0]   content_35;
  wire       [63:0]   content_36;
  wire       [63:0]   content_37;
  wire       [63:0]   content_38;
  wire       [63:0]   content_39;
  wire       [63:0]   content_40;
  wire       [63:0]   content_41;
  wire       [63:0]   content_42;
  wire       [63:0]   content_43;
  wire       [63:0]   content_44;
  wire       [63:0]   content_45;
  wire       [63:0]   content_46;
  wire       [63:0]   content_47;
  wire       [63:0]   content_48;
  wire       [63:0]   content_49;
  wire       [63:0]   content_50;
  wire       [63:0]   content_51;
  wire       [63:0]   content_52;
  wire       [63:0]   content_53;
  wire       [63:0]   content_54;
  wire       [63:0]   content_55;
  wire       [63:0]   content_56;
  wire       [63:0]   content_57;
  wire       [63:0]   content_58;
  wire       [63:0]   content_59;
  wire       [63:0]   content_60;
  wire       [63:0]   content_61;
  wire       [63:0]   content_62;
  wire       [63:0]   content_63;
  wire       [63:0]   content_64;
  wire       [63:0]   content_65;
  wire       [63:0]   content_66;
  wire       [63:0]   content_67;
  wire       [63:0]   content_68;
  wire       [63:0]   content_69;
  wire       [63:0]   content_70;
  wire       [63:0]   content_71;
  wire       [63:0]   content_72;
  wire       [63:0]   content_73;
  wire       [63:0]   content_74;
  wire       [63:0]   content_75;
  wire       [63:0]   content_76;
  wire       [63:0]   content_77;
  wire       [63:0]   content_78;
  wire       [63:0]   content_79;
  wire       [63:0]   content_80;
  wire       [63:0]   content_81;
  wire       [63:0]   content_82;
  wire       [63:0]   content_83;
  wire       [63:0]   content_84;
  wire       [63:0]   content_85;
  wire       [63:0]   content_86;
  wire       [63:0]   content_87;
  wire       [63:0]   content_88;
  wire       [63:0]   content_89;
  wire       [63:0]   content_90;
  wire       [63:0]   content_91;
  wire       [63:0]   content_92;
  wire       [63:0]   content_93;
  wire       [63:0]   content_94;
  wire       [63:0]   content_95;
  wire       [63:0]   content_96;
  wire       [63:0]   content_97;
  wire       [63:0]   content_98;
  wire       [63:0]   content_99;
  wire       [63:0]   content_100;
  wire       [63:0]   content_101;
  wire       [63:0]   content_102;
  wire       [63:0]   content_103;
  wire       [63:0]   content_104;
  wire       [63:0]   content_105;
  wire       [63:0]   content_106;
  wire       [63:0]   content_107;
  wire       [63:0]   content_108;
  wire       [63:0]   content_109;
  wire       [63:0]   content_110;
  wire       [63:0]   content_111;
  wire       [63:0]   content_112;
  wire       [63:0]   content_113;
  wire       [63:0]   content_114;
  wire       [63:0]   content_115;
  wire       [63:0]   content_116;
  wire       [63:0]   content_117;
  wire       [63:0]   content_118;
  wire       [63:0]   content_119;
  wire       [63:0]   content_120;
  wire       [63:0]   content_121;
  wire       [63:0]   content_122;
  wire       [63:0]   content_123;
  wire       [63:0]   content_124;
  wire       [63:0]   content_125;
  wire       [63:0]   content_126;
  wire       [63:0]   content_127;
  wire       [63:0]   content_128;
  wire       [63:0]   content_129;
  wire       [63:0]   content_130;
  wire       [63:0]   content_131;
  wire       [63:0]   content_132;
  wire       [63:0]   content_133;
  wire       [63:0]   content_134;
  wire       [63:0]   content_135;
  wire       [63:0]   content_136;
  wire       [63:0]   content_137;
  wire       [63:0]   content_138;
  wire       [63:0]   content_139;
  wire       [63:0]   content_140;
  wire       [63:0]   content_141;
  wire       [63:0]   content_142;
  wire       [63:0]   content_143;
  wire       [63:0]   content_144;
  wire       [63:0]   content_145;
  wire       [63:0]   content_146;
  wire       [63:0]   content_147;
  wire       [63:0]   content_148;
  wire       [63:0]   content_149;
  wire       [63:0]   content_150;
  wire       [63:0]   content_151;
  wire       [63:0]   content_152;
  wire       [63:0]   content_153;
  wire       [63:0]   content_154;
  wire       [63:0]   content_155;
  wire       [63:0]   content_156;
  wire       [63:0]   content_157;
  wire       [63:0]   content_158;
  wire       [63:0]   content_159;
  wire       [63:0]   content_160;
  wire       [63:0]   content_161;
  wire       [63:0]   content_162;
  wire       [63:0]   content_163;
  wire       [63:0]   content_164;
  wire       [63:0]   content_165;
  wire       [63:0]   content_166;
  wire       [63:0]   content_167;
  wire       [63:0]   content_168;
  wire       [63:0]   content_169;
  wire       [63:0]   content_170;
  wire       [63:0]   content_171;
  wire       [63:0]   content_172;
  wire       [63:0]   content_173;
  wire       [63:0]   content_174;
  wire       [63:0]   content_175;
  wire       [63:0]   content_176;
  wire       [63:0]   content_177;
  wire       [63:0]   content_178;
  wire       [63:0]   content_179;
  wire       [63:0]   content_180;
  wire       [63:0]   content_181;
  wire       [63:0]   content_182;
  wire       [63:0]   content_183;
  wire       [63:0]   content_184;
  wire       [63:0]   content_185;
  wire       [63:0]   content_186;
  wire       [63:0]   content_187;
  wire       [63:0]   content_188;
  wire       [63:0]   content_189;
  wire       [63:0]   content_190;
  wire       [63:0]   content_191;
  wire       [63:0]   content_192;
  wire       [63:0]   content_193;
  wire       [63:0]   content_194;
  wire       [63:0]   content_195;
  wire       [63:0]   content_196;
  wire       [63:0]   content_197;
  wire       [63:0]   content_198;
  wire       [63:0]   content_199;
  wire       [63:0]   content_200;
  wire       [63:0]   content_201;
  wire       [63:0]   content_202;
  wire       [63:0]   content_203;
  wire       [63:0]   content_204;
  wire       [63:0]   content_205;
  wire       [63:0]   content_206;
  wire       [63:0]   content_207;
  wire       [63:0]   content_208;
  wire       [63:0]   content_209;
  wire       [63:0]   content_210;
  wire       [63:0]   content_211;
  wire       [63:0]   content_212;
  wire       [63:0]   content_213;
  wire       [63:0]   content_214;
  wire       [63:0]   content_215;
  wire       [63:0]   content_216;
  wire       [63:0]   content_217;
  wire       [63:0]   content_218;
  wire       [63:0]   content_219;
  wire       [63:0]   content_220;
  wire       [63:0]   content_221;
  wire       [63:0]   content_222;
  wire       [63:0]   content_223;
  wire       [63:0]   content_224;
  wire       [63:0]   content_225;
  wire       [63:0]   content_226;
  wire       [63:0]   content_227;
  wire       [63:0]   content_228;
  wire       [63:0]   content_229;
  wire       [63:0]   content_230;
  wire       [63:0]   content_231;
  wire       [63:0]   content_232;
  wire       [63:0]   content_233;
  wire       [63:0]   content_234;
  wire       [63:0]   content_235;
  wire       [63:0]   content_236;
  wire       [63:0]   content_237;
  wire       [63:0]   content_238;
  wire       [63:0]   content_239;
  wire       [63:0]   content_240;
  wire       [63:0]   content_241;
  wire       [63:0]   content_242;
  wire       [63:0]   content_243;
  wire       [63:0]   content_244;
  wire       [63:0]   content_245;
  wire       [63:0]   content_246;
  wire       [63:0]   content_247;
  wire       [63:0]   content_248;
  wire       [63:0]   content_249;
  wire       [63:0]   content_250;
  wire       [63:0]   content_251;
  wire       [63:0]   content_252;
  wire       [63:0]   content_253;
  wire       [63:0]   content_254;
  wire       [63:0]   content_255;
  wire       [63:0]   content_256;
  wire       [63:0]   content_257;
  wire       [63:0]   content_258;
  wire       [63:0]   content_259;
  wire       [63:0]   content_260;
  wire       [63:0]   content_261;
  wire       [63:0]   content_262;
  wire       [63:0]   content_263;
  wire       [63:0]   content_264;
  wire       [63:0]   content_265;
  wire       [63:0]   content_266;
  wire       [63:0]   content_267;
  wire       [63:0]   content_268;
  wire       [63:0]   content_269;
  wire       [63:0]   content_270;
  wire       [63:0]   content_271;
  wire       [63:0]   content_272;
  wire       [63:0]   content_273;
  wire       [63:0]   content_274;
  wire       [63:0]   content_275;
  wire       [63:0]   content_276;
  wire       [63:0]   content_277;
  wire       [63:0]   content_278;
  wire       [63:0]   content_279;
  wire       [63:0]   content_280;
  wire       [63:0]   content_281;
  wire       [63:0]   content_282;
  wire       [63:0]   content_283;
  wire       [63:0]   content_284;
  wire       [63:0]   content_285;
  wire       [63:0]   content_286;
  wire       [63:0]   content_287;
  wire       [63:0]   content_288;
  wire       [63:0]   content_289;
  wire       [63:0]   content_290;
  wire       [63:0]   content_291;
  wire       [63:0]   content_292;
  wire       [63:0]   content_293;
  wire       [63:0]   content_294;
  wire       [63:0]   content_295;
  wire       [63:0]   content_296;
  wire       [63:0]   content_297;
  wire       [63:0]   content_298;
  wire       [63:0]   content_299;
  wire       [63:0]   content_300;
  wire       [63:0]   content_301;
  wire       [63:0]   content_302;
  wire       [63:0]   content_303;
  wire       [63:0]   content_304;
  wire       [63:0]   content_305;
  wire       [63:0]   content_306;
  wire       [63:0]   content_307;
  wire       [63:0]   content_308;
  wire       [63:0]   content_309;
  wire       [63:0]   content_310;
  wire       [63:0]   content_311;
  wire       [63:0]   content_312;
  wire       [63:0]   content_313;
  wire       [63:0]   content_314;
  wire       [63:0]   content_315;
  wire       [63:0]   content_316;
  wire       [63:0]   content_317;
  wire       [63:0]   content_318;
  wire       [63:0]   content_319;
  wire       [63:0]   content_320;
  wire       [63:0]   content_321;
  wire       [63:0]   content_322;
  wire       [63:0]   content_323;
  wire       [63:0]   content_324;
  wire       [63:0]   content_325;
  wire       [63:0]   content_326;
  wire       [63:0]   content_327;
  wire       [63:0]   content_328;
  wire       [63:0]   content_329;
  wire       [63:0]   content_330;
  wire       [63:0]   content_331;
  wire       [63:0]   content_332;
  wire       [63:0]   content_333;
  wire       [63:0]   content_334;
  wire       [63:0]   content_335;
  wire       [63:0]   content_336;
  wire       [63:0]   content_337;
  wire       [63:0]   content_338;
  wire       [63:0]   content_339;
  wire       [63:0]   content_340;
  wire       [63:0]   content_341;
  wire       [63:0]   content_342;
  wire       [63:0]   content_343;
  wire       [63:0]   content_344;
  wire       [63:0]   content_345;
  wire       [63:0]   content_346;
  wire       [63:0]   content_347;
  wire       [63:0]   content_348;
  wire       [63:0]   content_349;
  wire       [63:0]   content_350;
  wire       [63:0]   content_351;
  wire       [63:0]   content_352;
  wire       [63:0]   content_353;
  wire       [63:0]   content_354;
  wire       [63:0]   content_355;
  wire       [63:0]   content_356;
  wire       [63:0]   content_357;
  wire       [63:0]   content_358;
  wire       [63:0]   content_359;
  wire       [63:0]   content_360;
  wire       [63:0]   content_361;
  wire       [63:0]   content_362;
  wire       [63:0]   content_363;
  wire       [63:0]   content_364;
  wire       [63:0]   content_365;
  wire       [63:0]   content_366;
  wire       [63:0]   content_367;
  wire       [63:0]   content_368;
  wire       [63:0]   content_369;
  wire       [63:0]   content_370;
  wire       [63:0]   content_371;
  wire       [63:0]   content_372;
  wire       [63:0]   content_373;
  wire       [63:0]   content_374;
  wire       [63:0]   content_375;
  wire       [63:0]   content_376;
  wire       [63:0]   content_377;
  wire       [63:0]   content_378;
  wire       [63:0]   content_379;
  wire       [63:0]   content_380;
  wire       [63:0]   content_381;
  wire       [63:0]   content_382;
  wire       [63:0]   content_383;
  wire       [63:0]   content_384;
  wire       [63:0]   content_385;
  wire       [63:0]   content_386;
  wire       [63:0]   content_387;
  wire       [63:0]   content_388;
  wire       [63:0]   content_389;
  wire       [63:0]   content_390;
  wire       [63:0]   content_391;
  wire       [63:0]   content_392;
  wire       [63:0]   content_393;
  wire       [63:0]   content_394;
  wire       [63:0]   content_395;
  wire       [63:0]   content_396;
  wire       [63:0]   content_397;
  wire       [63:0]   content_398;
  wire       [63:0]   content_399;
  wire       [63:0]   content_400;
  wire       [63:0]   content_401;
  wire       [63:0]   content_402;
  wire       [63:0]   content_403;
  wire       [63:0]   content_404;
  wire       [63:0]   content_405;
  wire       [63:0]   content_406;
  wire       [63:0]   content_407;
  wire       [63:0]   content_408;
  wire       [63:0]   content_409;
  wire       [63:0]   content_410;
  wire       [63:0]   content_411;
  wire       [63:0]   content_412;
  wire       [63:0]   content_413;
  wire       [63:0]   content_414;
  wire       [63:0]   content_415;
  wire       [63:0]   content_416;
  wire       [63:0]   content_417;
  wire       [63:0]   content_418;
  wire       [63:0]   content_419;
  wire       [63:0]   content_420;
  wire       [63:0]   content_421;
  wire       [63:0]   content_422;
  wire       [63:0]   content_423;
  wire       [63:0]   content_424;
  wire       [63:0]   content_425;
  wire       [63:0]   content_426;
  wire       [63:0]   content_427;
  wire       [63:0]   content_428;
  wire       [63:0]   content_429;
  wire       [63:0]   content_430;
  wire       [63:0]   content_431;
  wire       [63:0]   content_432;
  wire       [63:0]   content_433;
  wire       [63:0]   content_434;
  wire       [63:0]   content_435;
  wire       [63:0]   content_436;
  wire       [63:0]   content_437;
  wire       [63:0]   content_438;
  wire       [63:0]   content_439;
  wire       [63:0]   content_440;
  wire       [63:0]   content_441;
  wire       [63:0]   content_442;
  wire       [63:0]   content_443;
  wire       [63:0]   content_444;
  wire       [63:0]   content_445;
  wire       [63:0]   content_446;
  wire       [63:0]   content_447;
  wire       [63:0]   content_448;
  wire       [63:0]   content_449;
  wire       [63:0]   content_450;
  wire       [63:0]   content_451;
  wire       [63:0]   content_452;
  wire       [63:0]   content_453;
  wire       [63:0]   content_454;
  wire       [63:0]   content_455;
  wire       [63:0]   content_456;
  wire       [63:0]   content_457;
  wire       [63:0]   content_458;
  wire       [63:0]   content_459;
  wire       [63:0]   content_460;
  wire       [63:0]   content_461;
  wire       [63:0]   content_462;
  wire       [63:0]   content_463;
  wire       [63:0]   content_464;
  wire       [63:0]   content_465;
  wire       [63:0]   content_466;
  wire       [63:0]   content_467;
  wire       [63:0]   content_468;
  wire       [63:0]   content_469;
  wire       [63:0]   content_470;
  wire       [63:0]   content_471;
  wire       [63:0]   content_472;
  wire       [63:0]   content_473;
  wire       [63:0]   content_474;
  wire       [63:0]   content_475;
  wire       [63:0]   content_476;
  wire       [63:0]   content_477;
  wire       [63:0]   content_478;
  wire       [63:0]   content_479;
  wire       [63:0]   content_480;
  wire       [63:0]   content_481;
  wire       [63:0]   content_482;
  wire       [63:0]   content_483;
  wire       [63:0]   content_484;
  wire       [63:0]   content_485;
  wire       [63:0]   content_486;
  wire       [63:0]   content_487;
  wire       [63:0]   content_488;
  wire       [63:0]   content_489;
  wire       [63:0]   content_490;
  wire       [63:0]   content_491;
  wire       [63:0]   content_492;
  wire       [63:0]   content_493;
  wire       [63:0]   content_494;
  wire       [63:0]   content_495;
  wire       [63:0]   content_496;
  wire       [63:0]   content_497;
  wire       [63:0]   content_498;
  wire       [63:0]   content_499;
  wire       [63:0]   content_500;
  wire       [63:0]   content_501;
  wire       [63:0]   content_502;
  wire       [63:0]   content_503;
  wire       [63:0]   content_504;
  wire       [63:0]   content_505;
  wire       [63:0]   content_506;
  wire       [63:0]   content_507;
  wire       [63:0]   content_508;
  wire       [63:0]   content_509;
  wire       [63:0]   content_510;
  wire       [63:0]   content_511;
  wire       [63:0]   content_512;
  wire       [63:0]   content_513;
  wire       [63:0]   content_514;
  wire       [63:0]   content_515;
  wire       [63:0]   content_516;
  wire       [63:0]   content_517;
  wire       [63:0]   content_518;
  wire       [63:0]   content_519;
  wire       [63:0]   content_520;
  wire       [63:0]   content_521;
  wire       [63:0]   content_522;
  wire       [63:0]   content_523;
  wire       [63:0]   content_524;
  wire       [63:0]   content_525;
  wire       [63:0]   content_526;
  wire       [63:0]   content_527;
  wire       [63:0]   content_528;
  wire       [63:0]   content_529;
  wire       [63:0]   content_530;
  wire       [63:0]   content_531;
  wire       [63:0]   content_532;
  wire       [63:0]   content_533;
  wire       [63:0]   content_534;
  wire       [63:0]   content_535;
  wire       [63:0]   content_536;
  wire       [63:0]   content_537;
  wire       [63:0]   content_538;
  wire       [63:0]   content_539;
  wire       [63:0]   content_540;
  wire       [63:0]   content_541;
  wire       [63:0]   content_542;
  wire       [63:0]   content_543;
  wire       [63:0]   content_544;
  wire       [63:0]   content_545;
  wire       [63:0]   content_546;
  wire       [63:0]   content_547;
  wire       [63:0]   content_548;
  wire       [63:0]   content_549;
  wire       [63:0]   content_550;
  wire       [63:0]   content_551;
  wire       [63:0]   content_552;
  wire       [63:0]   content_553;
  wire       [63:0]   content_554;
  wire       [63:0]   content_555;
  wire       [63:0]   content_556;
  wire       [63:0]   content_557;
  wire       [63:0]   content_558;
  wire       [63:0]   content_559;
  wire       [63:0]   content_560;
  wire       [63:0]   content_561;
  wire       [63:0]   content_562;
  wire       [63:0]   content_563;
  wire       [63:0]   content_564;
  wire       [63:0]   content_565;
  wire       [63:0]   content_566;
  wire       [63:0]   content_567;
  wire       [63:0]   content_568;
  wire       [63:0]   content_569;
  wire       [63:0]   content_570;
  wire       [63:0]   content_571;
  wire       [63:0]   content_572;
  wire       [63:0]   content_573;
  wire       [63:0]   content_574;
  wire       [63:0]   content_575;
  wire       [63:0]   content_576;
  wire       [63:0]   content_577;
  wire       [63:0]   content_578;
  wire       [63:0]   content_579;
  wire       [63:0]   content_580;
  wire       [63:0]   content_581;
  wire       [63:0]   content_582;
  wire       [63:0]   content_583;
  wire       [63:0]   content_584;
  wire       [63:0]   content_585;
  wire       [63:0]   content_586;
  wire       [63:0]   content_587;
  wire       [63:0]   content_588;
  wire       [63:0]   content_589;
  wire       [63:0]   content_590;
  wire       [63:0]   content_591;
  wire       [63:0]   content_592;
  wire       [63:0]   content_593;
  wire       [63:0]   content_594;
  wire       [63:0]   content_595;
  wire       [63:0]   content_596;
  wire       [63:0]   content_597;
  wire       [63:0]   content_598;
  wire       [63:0]   content_599;
  wire       [63:0]   content_600;
  wire       [63:0]   content_601;
  wire       [63:0]   content_602;
  wire       [63:0]   content_603;
  wire       [63:0]   content_604;
  wire       [63:0]   content_605;
  wire       [63:0]   content_606;
  wire       [63:0]   content_607;
  wire       [63:0]   content_608;
  wire       [63:0]   content_609;
  wire       [63:0]   content_610;
  wire       [63:0]   content_611;
  wire       [63:0]   content_612;
  wire       [63:0]   content_613;
  wire       [63:0]   content_614;
  wire       [63:0]   content_615;
  wire       [63:0]   content_616;
  wire       [63:0]   content_617;
  wire       [63:0]   content_618;
  wire       [63:0]   content_619;
  wire       [63:0]   content_620;
  wire       [63:0]   content_621;
  wire       [63:0]   content_622;
  wire       [63:0]   content_623;
  wire       [63:0]   content_624;
  wire       [63:0]   content_625;
  wire       [63:0]   content_626;
  wire       [63:0]   content_627;
  wire       [63:0]   content_628;
  wire       [63:0]   content_629;
  wire       [63:0]   content_630;
  wire       [63:0]   content_631;
  wire       [63:0]   content_632;
  wire       [63:0]   content_633;
  wire       [63:0]   content_634;
  wire       [63:0]   content_635;
  wire       [63:0]   content_636;
  wire       [63:0]   content_637;
  wire       [63:0]   content_638;
  wire       [63:0]   content_639;
  wire       [63:0]   content_640;
  wire       [63:0]   content_641;
  wire       [63:0]   content_642;
  wire       [63:0]   content_643;
  wire       [63:0]   content_644;
  wire       [63:0]   content_645;
  wire       [63:0]   content_646;
  wire       [63:0]   content_647;
  wire       [63:0]   content_648;
  wire       [63:0]   content_649;
  wire       [63:0]   content_650;
  wire       [63:0]   content_651;
  wire       [63:0]   content_652;
  wire       [63:0]   content_653;
  wire       [63:0]   content_654;
  wire       [63:0]   content_655;
  wire       [63:0]   content_656;
  wire       [63:0]   content_657;
  wire       [63:0]   content_658;
  wire       [63:0]   content_659;
  wire       [63:0]   content_660;
  wire       [63:0]   content_661;
  wire       [63:0]   content_662;
  wire       [63:0]   content_663;
  wire       [63:0]   content_664;
  wire       [63:0]   content_665;
  wire       [63:0]   content_666;
  wire       [63:0]   content_667;
  wire       [63:0]   content_668;
  wire       [63:0]   content_669;
  wire       [63:0]   content_670;
  wire       [63:0]   content_671;
  wire       [63:0]   content_672;
  wire       [63:0]   content_673;
  wire       [63:0]   content_674;
  wire       [63:0]   content_675;
  wire       [63:0]   content_676;
  wire       [63:0]   content_677;
  wire       [63:0]   content_678;
  wire       [63:0]   content_679;
  wire       [63:0]   content_680;
  wire       [63:0]   content_681;
  wire       [63:0]   content_682;
  wire       [63:0]   content_683;
  wire       [63:0]   content_684;
  wire       [63:0]   content_685;
  wire       [63:0]   content_686;
  wire       [63:0]   content_687;
  wire       [63:0]   content_688;
  wire       [63:0]   content_689;
  wire       [63:0]   content_690;
  wire       [63:0]   content_691;
  wire       [63:0]   content_692;
  wire       [63:0]   content_693;
  wire       [63:0]   content_694;
  wire       [63:0]   content_695;
  wire       [63:0]   content_696;
  wire       [63:0]   content_697;
  wire       [63:0]   content_698;
  wire       [63:0]   content_699;
  wire       [63:0]   content_700;
  wire       [63:0]   content_701;
  wire       [63:0]   content_702;
  wire       [63:0]   content_703;
  wire       [63:0]   content_704;
  wire       [63:0]   content_705;
  wire       [63:0]   content_706;
  wire       [63:0]   content_707;
  wire       [63:0]   content_708;
  wire       [63:0]   content_709;
  wire       [63:0]   content_710;
  wire       [63:0]   content_711;
  wire       [63:0]   content_712;
  wire       [63:0]   content_713;
  wire       [63:0]   content_714;
  wire       [63:0]   content_715;
  wire       [63:0]   content_716;
  wire       [63:0]   content_717;
  wire       [63:0]   content_718;
  wire       [63:0]   content_719;
  wire       [63:0]   content_720;
  wire       [63:0]   content_721;
  wire       [63:0]   content_722;
  wire       [63:0]   content_723;
  wire       [63:0]   content_724;
  wire       [63:0]   content_725;
  wire       [63:0]   content_726;
  wire       [63:0]   content_727;
  wire       [63:0]   content_728;
  wire       [63:0]   content_729;
  wire       [63:0]   content_730;
  wire       [63:0]   content_731;
  wire       [63:0]   content_732;
  wire       [63:0]   content_733;
  wire       [63:0]   content_734;
  wire       [63:0]   content_735;
  wire       [63:0]   content_736;
  wire       [63:0]   content_737;
  wire       [63:0]   content_738;
  wire       [63:0]   content_739;
  wire       [63:0]   content_740;
  wire       [63:0]   content_741;
  wire       [63:0]   content_742;
  wire       [63:0]   content_743;
  wire       [63:0]   content_744;
  wire       [63:0]   content_745;
  wire       [63:0]   content_746;
  wire       [63:0]   content_747;
  wire       [63:0]   content_748;
  wire       [63:0]   content_749;
  wire       [63:0]   content_750;
  wire       [63:0]   content_751;
  wire       [63:0]   content_752;
  wire       [63:0]   content_753;
  wire       [63:0]   content_754;
  wire       [63:0]   content_755;
  wire       [63:0]   content_756;
  wire       [63:0]   content_757;
  wire       [63:0]   content_758;
  wire       [63:0]   content_759;
  wire       [63:0]   content_760;
  wire       [63:0]   content_761;
  wire       [63:0]   content_762;
  wire       [63:0]   content_763;
  wire       [63:0]   content_764;
  wire       [63:0]   content_765;
  wire       [63:0]   content_766;
  wire       [63:0]   content_767;
  wire       [63:0]   content_768;
  wire       [63:0]   content_769;
  wire       [63:0]   content_770;
  wire       [63:0]   content_771;
  wire       [63:0]   content_772;
  wire       [63:0]   content_773;
  wire       [63:0]   content_774;
  wire       [63:0]   content_775;
  wire       [63:0]   content_776;
  wire       [63:0]   content_777;
  wire       [63:0]   content_778;
  wire       [63:0]   content_779;
  wire       [63:0]   content_780;
  wire       [63:0]   content_781;
  wire       [63:0]   content_782;
  wire       [63:0]   content_783;
  wire       [63:0]   content_784;
  wire       [63:0]   content_785;
  wire       [63:0]   content_786;
  wire       [63:0]   content_787;
  wire       [63:0]   content_788;
  wire       [63:0]   content_789;
  wire       [63:0]   content_790;
  wire       [63:0]   content_791;
  wire       [63:0]   content_792;
  wire       [63:0]   content_793;
  wire       [63:0]   content_794;
  wire       [63:0]   content_795;
  wire       [63:0]   content_796;
  wire       [63:0]   content_797;
  wire       [63:0]   content_798;
  wire       [63:0]   content_799;
  wire       [63:0]   content_800;
  wire       [63:0]   content_801;
  wire       [63:0]   content_802;
  wire       [63:0]   content_803;
  wire       [63:0]   content_804;
  wire       [63:0]   content_805;
  wire       [63:0]   content_806;
  wire       [63:0]   content_807;
  wire       [63:0]   content_808;
  wire       [63:0]   content_809;
  wire       [63:0]   content_810;
  wire       [63:0]   content_811;
  wire       [63:0]   content_812;
  wire       [63:0]   content_813;
  wire       [63:0]   content_814;
  wire       [63:0]   content_815;
  wire       [63:0]   content_816;
  wire       [63:0]   content_817;
  wire       [63:0]   content_818;
  wire       [63:0]   content_819;
  wire       [63:0]   content_820;
  wire       [63:0]   content_821;
  wire       [63:0]   content_822;
  wire       [63:0]   content_823;
  wire       [63:0]   content_824;
  wire       [63:0]   content_825;
  wire       [63:0]   content_826;
  wire       [63:0]   content_827;
  wire       [63:0]   content_828;
  wire       [63:0]   content_829;
  wire       [63:0]   content_830;
  wire       [63:0]   content_831;
  wire       [63:0]   content_832;
  wire       [63:0]   content_833;
  wire       [63:0]   content_834;
  wire       [63:0]   content_835;
  wire       [63:0]   content_836;
  wire       [63:0]   content_837;
  wire       [63:0]   content_838;
  wire       [63:0]   content_839;
  wire       [63:0]   content_840;
  wire       [63:0]   content_841;
  wire       [63:0]   content_842;
  wire       [63:0]   content_843;
  wire       [63:0]   content_844;
  wire       [63:0]   content_845;
  wire       [63:0]   content_846;
  wire       [63:0]   content_847;
  wire       [63:0]   content_848;
  wire       [63:0]   content_849;
  wire       [63:0]   content_850;
  wire       [63:0]   content_851;
  wire       [63:0]   content_852;
  wire       [63:0]   content_853;
  wire       [63:0]   content_854;
  wire       [63:0]   content_855;
  wire       [63:0]   content_856;
  wire       [63:0]   content_857;
  wire       [63:0]   content_858;
  wire       [63:0]   content_859;
  wire       [63:0]   content_860;
  wire       [63:0]   content_861;
  wire       [63:0]   content_862;
  wire       [63:0]   content_863;
  wire       [63:0]   content_864;
  wire       [63:0]   content_865;
  wire       [63:0]   content_866;
  wire       [63:0]   content_867;
  wire       [63:0]   content_868;
  wire       [63:0]   content_869;
  wire       [63:0]   content_870;
  wire       [63:0]   content_871;
  wire       [63:0]   content_872;
  wire       [63:0]   content_873;
  wire       [63:0]   content_874;
  wire       [63:0]   content_875;
  wire       [63:0]   content_876;
  wire       [63:0]   content_877;
  wire       [63:0]   content_878;
  wire       [63:0]   content_879;
  wire       [63:0]   content_880;
  wire       [63:0]   content_881;
  wire       [63:0]   content_882;
  wire       [63:0]   content_883;
  wire       [63:0]   content_884;
  wire       [63:0]   content_885;
  wire       [63:0]   content_886;
  wire       [63:0]   content_887;
  wire       [63:0]   content_888;
  wire       [63:0]   content_889;
  wire       [63:0]   content_890;
  wire       [63:0]   content_891;
  wire       [63:0]   content_892;
  wire       [63:0]   content_893;
  wire       [63:0]   content_894;
  wire       [63:0]   content_895;
  wire       [63:0]   content_896;
  wire       [63:0]   content_897;
  wire       [63:0]   content_898;
  wire       [63:0]   content_899;
  wire       [63:0]   content_900;
  wire       [63:0]   content_901;
  wire       [63:0]   content_902;
  wire       [63:0]   content_903;
  wire       [63:0]   content_904;
  wire       [63:0]   content_905;
  wire       [63:0]   content_906;
  wire       [63:0]   content_907;
  wire       [63:0]   content_908;
  wire       [63:0]   content_909;
  wire       [63:0]   content_910;
  wire       [63:0]   content_911;
  wire       [63:0]   content_912;
  wire       [63:0]   content_913;
  wire       [63:0]   content_914;
  wire       [63:0]   content_915;
  wire       [63:0]   content_916;
  wire       [63:0]   content_917;
  wire       [63:0]   content_918;
  wire       [63:0]   content_919;
  wire       [63:0]   content_920;
  wire       [63:0]   content_921;
  wire       [63:0]   content_922;
  wire       [63:0]   content_923;
  wire       [63:0]   content_924;
  wire       [63:0]   content_925;
  wire       [63:0]   content_926;
  wire       [63:0]   content_927;
  wire       [63:0]   content_928;
  wire       [63:0]   content_929;
  wire       [63:0]   content_930;
  wire       [63:0]   content_931;
  wire       [63:0]   content_932;
  wire       [63:0]   content_933;
  wire       [63:0]   content_934;
  wire       [63:0]   content_935;
  wire       [63:0]   content_936;
  wire       [63:0]   content_937;
  wire       [63:0]   content_938;
  wire       [63:0]   content_939;
  wire       [63:0]   content_940;
  wire       [63:0]   content_941;
  wire       [63:0]   content_942;
  wire       [63:0]   content_943;
  wire       [63:0]   content_944;
  wire       [63:0]   content_945;
  wire       [63:0]   content_946;
  wire       [63:0]   content_947;
  wire       [63:0]   content_948;
  wire       [63:0]   content_949;
  wire       [63:0]   content_950;
  wire       [63:0]   content_951;
  wire       [63:0]   content_952;
  wire       [63:0]   content_953;
  wire       [63:0]   content_954;
  wire       [63:0]   content_955;
  wire       [63:0]   content_956;
  wire       [63:0]   content_957;
  wire       [63:0]   content_958;
  wire       [63:0]   content_959;
  wire       [63:0]   content_960;
  wire       [63:0]   content_961;
  wire       [63:0]   content_962;
  wire       [63:0]   content_963;
  wire       [63:0]   content_964;
  wire       [63:0]   content_965;
  wire       [63:0]   content_966;
  wire       [63:0]   content_967;
  wire       [63:0]   content_968;
  wire       [63:0]   content_969;
  wire       [63:0]   content_970;
  wire       [63:0]   content_971;
  wire       [63:0]   content_972;
  wire       [63:0]   content_973;
  wire       [63:0]   content_974;
  wire       [63:0]   content_975;
  wire       [63:0]   content_976;
  wire       [63:0]   content_977;
  wire       [63:0]   content_978;
  wire       [63:0]   content_979;
  wire       [63:0]   content_980;
  wire       [63:0]   content_981;
  wire       [63:0]   content_982;
  wire       [63:0]   content_983;
  wire       [63:0]   content_984;
  wire       [63:0]   content_985;
  wire       [63:0]   content_986;
  wire       [63:0]   content_987;
  wire       [63:0]   content_988;
  wire       [63:0]   content_989;
  wire       [63:0]   content_990;
  wire       [63:0]   content_991;
  wire       [63:0]   content_992;
  wire       [63:0]   content_993;
  wire       [63:0]   content_994;
  wire       [63:0]   content_995;
  wire       [63:0]   content_996;
  wire       [63:0]   content_997;
  wire       [63:0]   content_998;
  wire       [63:0]   content_999;
  wire       [63:0]   content_1000;
  wire       [63:0]   content_1001;
  wire       [63:0]   content_1002;
  wire       [63:0]   content_1003;
  wire       [63:0]   content_1004;
  wire       [63:0]   content_1005;
  wire       [63:0]   content_1006;
  wire       [63:0]   content_1007;
  wire       [63:0]   content_1008;
  wire       [63:0]   content_1009;
  wire       [63:0]   content_1010;
  wire       [63:0]   content_1011;
  wire       [63:0]   content_1012;
  wire       [63:0]   content_1013;
  wire       [63:0]   content_1014;
  wire       [63:0]   content_1015;
  wire       [63:0]   content_1016;
  wire       [63:0]   content_1017;
  wire       [63:0]   content_1018;
  wire       [63:0]   content_1019;
  wire       [63:0]   content_1020;
  wire       [63:0]   content_1021;
  wire       [63:0]   content_1022;
  wire       [63:0]   content_1023;
  wire       [9:0]    _zz_1_;
  reg [63:0] mem [0:1023];

  assign _zz_3_ = (address >>> 3);
  initial begin
    $readmemb("dataMem.v_toplevel_mem.bin",mem);
  end
  assign _zz_2_ = mem[_zz_1_];
  always @ (posedge clk) begin
    if(memWrite) begin
      mem[_zz_3_] <= writeData;
    end
  end

  assign content_0 = 64'h0;
  assign content_1 = 64'h0000000000000001;
  assign content_2 = 64'h0000000000000002;
  assign content_3 = 64'h0000000000000003;
  assign content_4 = 64'h0000000000000004;
  assign content_5 = 64'h0000000000000005;
  assign content_6 = 64'h0000000000000006;
  assign content_7 = 64'h0000000000000007;
  assign content_8 = 64'h0000000000000008;
  assign content_9 = 64'h0000000000000009;
  assign content_10 = 64'h000000000000000a;
  assign content_11 = 64'h000000000000000b;
  assign content_12 = 64'h000000000000000c;
  assign content_13 = 64'h000000000000000d;
  assign content_14 = 64'h000000000000000e;
  assign content_15 = 64'h000000000000000f;
  assign content_16 = 64'h0000000000000010;
  assign content_17 = 64'h0000000000000011;
  assign content_18 = 64'h0000000000000012;
  assign content_19 = 64'h0000000000000013;
  assign content_20 = 64'h0000000000000014;
  assign content_21 = 64'h0000000000000015;
  assign content_22 = 64'h0000000000000016;
  assign content_23 = 64'h0000000000000017;
  assign content_24 = 64'h0000000000000018;
  assign content_25 = 64'h0000000000000019;
  assign content_26 = 64'h000000000000001a;
  assign content_27 = 64'h000000000000001b;
  assign content_28 = 64'h000000000000001c;
  assign content_29 = 64'h000000000000001d;
  assign content_30 = 64'h000000000000001e;
  assign content_31 = 64'h000000000000001f;
  assign content_32 = 64'h0000000000000020;
  assign content_33 = 64'h0000000000000021;
  assign content_34 = 64'h0000000000000022;
  assign content_35 = 64'h0000000000000023;
  assign content_36 = 64'h0000000000000024;
  assign content_37 = 64'h0000000000000025;
  assign content_38 = 64'h0000000000000026;
  assign content_39 = 64'h0000000000000027;
  assign content_40 = 64'h0000000000000028;
  assign content_41 = 64'h0000000000000029;
  assign content_42 = 64'h000000000000002a;
  assign content_43 = 64'h000000000000002b;
  assign content_44 = 64'h000000000000002c;
  assign content_45 = 64'h000000000000002d;
  assign content_46 = 64'h000000000000002e;
  assign content_47 = 64'h000000000000002f;
  assign content_48 = 64'h0000000000000030;
  assign content_49 = 64'h0000000000000031;
  assign content_50 = 64'h0000000000000032;
  assign content_51 = 64'h0000000000000033;
  assign content_52 = 64'h0000000000000034;
  assign content_53 = 64'h0000000000000035;
  assign content_54 = 64'h0000000000000036;
  assign content_55 = 64'h0000000000000037;
  assign content_56 = 64'h0000000000000038;
  assign content_57 = 64'h0000000000000039;
  assign content_58 = 64'h000000000000003a;
  assign content_59 = 64'h000000000000003b;
  assign content_60 = 64'h000000000000003c;
  assign content_61 = 64'h000000000000003d;
  assign content_62 = 64'h000000000000003e;
  assign content_63 = 64'h000000000000003f;
  assign content_64 = 64'h0000000000000040;
  assign content_65 = 64'h0000000000000041;
  assign content_66 = 64'h0000000000000042;
  assign content_67 = 64'h0000000000000043;
  assign content_68 = 64'h0000000000000044;
  assign content_69 = 64'h0000000000000045;
  assign content_70 = 64'h0000000000000046;
  assign content_71 = 64'h0000000000000047;
  assign content_72 = 64'h0000000000000048;
  assign content_73 = 64'h0000000000000049;
  assign content_74 = 64'h000000000000004a;
  assign content_75 = 64'h000000000000004b;
  assign content_76 = 64'h000000000000004c;
  assign content_77 = 64'h000000000000004d;
  assign content_78 = 64'h000000000000004e;
  assign content_79 = 64'h000000000000004f;
  assign content_80 = 64'h0000000000000050;
  assign content_81 = 64'h0000000000000051;
  assign content_82 = 64'h0000000000000052;
  assign content_83 = 64'h0000000000000053;
  assign content_84 = 64'h0000000000000054;
  assign content_85 = 64'h0000000000000055;
  assign content_86 = 64'h0000000000000056;
  assign content_87 = 64'h0000000000000057;
  assign content_88 = 64'h0000000000000058;
  assign content_89 = 64'h0000000000000059;
  assign content_90 = 64'h000000000000005a;
  assign content_91 = 64'h000000000000005b;
  assign content_92 = 64'h000000000000005c;
  assign content_93 = 64'h000000000000005d;
  assign content_94 = 64'h000000000000005e;
  assign content_95 = 64'h000000000000005f;
  assign content_96 = 64'h0000000000000060;
  assign content_97 = 64'h0000000000000061;
  assign content_98 = 64'h0000000000000062;
  assign content_99 = 64'h0000000000000063;
  assign content_100 = 64'h0000000000000064;
  assign content_101 = 64'h0000000000000065;
  assign content_102 = 64'h0000000000000066;
  assign content_103 = 64'h0000000000000067;
  assign content_104 = 64'h0000000000000068;
  assign content_105 = 64'h0000000000000069;
  assign content_106 = 64'h000000000000006a;
  assign content_107 = 64'h000000000000006b;
  assign content_108 = 64'h000000000000006c;
  assign content_109 = 64'h000000000000006d;
  assign content_110 = 64'h000000000000006e;
  assign content_111 = 64'h000000000000006f;
  assign content_112 = 64'h0000000000000070;
  assign content_113 = 64'h0000000000000071;
  assign content_114 = 64'h0000000000000072;
  assign content_115 = 64'h0000000000000073;
  assign content_116 = 64'h0000000000000074;
  assign content_117 = 64'h0000000000000075;
  assign content_118 = 64'h0000000000000076;
  assign content_119 = 64'h0000000000000077;
  assign content_120 = 64'h0000000000000078;
  assign content_121 = 64'h0000000000000079;
  assign content_122 = 64'h000000000000007a;
  assign content_123 = 64'h000000000000007b;
  assign content_124 = 64'h000000000000007c;
  assign content_125 = 64'h000000000000007d;
  assign content_126 = 64'h000000000000007e;
  assign content_127 = 64'h000000000000007f;
  assign content_128 = 64'h0000000000000080;
  assign content_129 = 64'h0000000000000081;
  assign content_130 = 64'h0000000000000082;
  assign content_131 = 64'h0000000000000083;
  assign content_132 = 64'h0000000000000084;
  assign content_133 = 64'h0000000000000085;
  assign content_134 = 64'h0000000000000086;
  assign content_135 = 64'h0000000000000087;
  assign content_136 = 64'h0000000000000088;
  assign content_137 = 64'h0000000000000089;
  assign content_138 = 64'h000000000000008a;
  assign content_139 = 64'h000000000000008b;
  assign content_140 = 64'h000000000000008c;
  assign content_141 = 64'h000000000000008d;
  assign content_142 = 64'h000000000000008e;
  assign content_143 = 64'h000000000000008f;
  assign content_144 = 64'h0000000000000090;
  assign content_145 = 64'h0000000000000091;
  assign content_146 = 64'h0000000000000092;
  assign content_147 = 64'h0000000000000093;
  assign content_148 = 64'h0000000000000094;
  assign content_149 = 64'h0000000000000095;
  assign content_150 = 64'h0000000000000096;
  assign content_151 = 64'h0000000000000097;
  assign content_152 = 64'h0000000000000098;
  assign content_153 = 64'h0000000000000099;
  assign content_154 = 64'h000000000000009a;
  assign content_155 = 64'h000000000000009b;
  assign content_156 = 64'h000000000000009c;
  assign content_157 = 64'h000000000000009d;
  assign content_158 = 64'h000000000000009e;
  assign content_159 = 64'h000000000000009f;
  assign content_160 = 64'h00000000000000a0;
  assign content_161 = 64'h00000000000000a1;
  assign content_162 = 64'h00000000000000a2;
  assign content_163 = 64'h00000000000000a3;
  assign content_164 = 64'h00000000000000a4;
  assign content_165 = 64'h00000000000000a5;
  assign content_166 = 64'h00000000000000a6;
  assign content_167 = 64'h00000000000000a7;
  assign content_168 = 64'h00000000000000a8;
  assign content_169 = 64'h00000000000000a9;
  assign content_170 = 64'h00000000000000aa;
  assign content_171 = 64'h00000000000000ab;
  assign content_172 = 64'h00000000000000ac;
  assign content_173 = 64'h00000000000000ad;
  assign content_174 = 64'h00000000000000ae;
  assign content_175 = 64'h00000000000000af;
  assign content_176 = 64'h00000000000000b0;
  assign content_177 = 64'h00000000000000b1;
  assign content_178 = 64'h00000000000000b2;
  assign content_179 = 64'h00000000000000b3;
  assign content_180 = 64'h00000000000000b4;
  assign content_181 = 64'h00000000000000b5;
  assign content_182 = 64'h00000000000000b6;
  assign content_183 = 64'h00000000000000b7;
  assign content_184 = 64'h00000000000000b8;
  assign content_185 = 64'h00000000000000b9;
  assign content_186 = 64'h00000000000000ba;
  assign content_187 = 64'h00000000000000bb;
  assign content_188 = 64'h00000000000000bc;
  assign content_189 = 64'h00000000000000bd;
  assign content_190 = 64'h00000000000000be;
  assign content_191 = 64'h00000000000000bf;
  assign content_192 = 64'h00000000000000c0;
  assign content_193 = 64'h00000000000000c1;
  assign content_194 = 64'h00000000000000c2;
  assign content_195 = 64'h00000000000000c3;
  assign content_196 = 64'h00000000000000c4;
  assign content_197 = 64'h00000000000000c5;
  assign content_198 = 64'h00000000000000c6;
  assign content_199 = 64'h00000000000000c7;
  assign content_200 = 64'h00000000000000c8;
  assign content_201 = 64'h00000000000000c9;
  assign content_202 = 64'h00000000000000ca;
  assign content_203 = 64'h00000000000000cb;
  assign content_204 = 64'h00000000000000cc;
  assign content_205 = 64'h00000000000000cd;
  assign content_206 = 64'h00000000000000ce;
  assign content_207 = 64'h00000000000000cf;
  assign content_208 = 64'h00000000000000d0;
  assign content_209 = 64'h00000000000000d1;
  assign content_210 = 64'h00000000000000d2;
  assign content_211 = 64'h00000000000000d3;
  assign content_212 = 64'h00000000000000d4;
  assign content_213 = 64'h00000000000000d5;
  assign content_214 = 64'h00000000000000d6;
  assign content_215 = 64'h00000000000000d7;
  assign content_216 = 64'h00000000000000d8;
  assign content_217 = 64'h00000000000000d9;
  assign content_218 = 64'h00000000000000da;
  assign content_219 = 64'h00000000000000db;
  assign content_220 = 64'h00000000000000dc;
  assign content_221 = 64'h00000000000000dd;
  assign content_222 = 64'h00000000000000de;
  assign content_223 = 64'h00000000000000df;
  assign content_224 = 64'h00000000000000e0;
  assign content_225 = 64'h00000000000000e1;
  assign content_226 = 64'h00000000000000e2;
  assign content_227 = 64'h00000000000000e3;
  assign content_228 = 64'h00000000000000e4;
  assign content_229 = 64'h00000000000000e5;
  assign content_230 = 64'h00000000000000e6;
  assign content_231 = 64'h00000000000000e7;
  assign content_232 = 64'h00000000000000e8;
  assign content_233 = 64'h00000000000000e9;
  assign content_234 = 64'h00000000000000ea;
  assign content_235 = 64'h00000000000000eb;
  assign content_236 = 64'h00000000000000ec;
  assign content_237 = 64'h00000000000000ed;
  assign content_238 = 64'h00000000000000ee;
  assign content_239 = 64'h00000000000000ef;
  assign content_240 = 64'h00000000000000f0;
  assign content_241 = 64'h00000000000000f1;
  assign content_242 = 64'h00000000000000f2;
  assign content_243 = 64'h00000000000000f3;
  assign content_244 = 64'h00000000000000f4;
  assign content_245 = 64'h00000000000000f5;
  assign content_246 = 64'h00000000000000f6;
  assign content_247 = 64'h00000000000000f7;
  assign content_248 = 64'h00000000000000f8;
  assign content_249 = 64'h00000000000000f9;
  assign content_250 = 64'h00000000000000fa;
  assign content_251 = 64'h00000000000000fb;
  assign content_252 = 64'h00000000000000fc;
  assign content_253 = 64'h00000000000000fd;
  assign content_254 = 64'h00000000000000fe;
  assign content_255 = 64'h00000000000000ff;
  assign content_256 = 64'h0000000000000100;
  assign content_257 = 64'h0000000000000101;
  assign content_258 = 64'h0000000000000102;
  assign content_259 = 64'h0000000000000103;
  assign content_260 = 64'h0000000000000104;
  assign content_261 = 64'h0000000000000105;
  assign content_262 = 64'h0000000000000106;
  assign content_263 = 64'h0000000000000107;
  assign content_264 = 64'h0000000000000108;
  assign content_265 = 64'h0000000000000109;
  assign content_266 = 64'h000000000000010a;
  assign content_267 = 64'h000000000000010b;
  assign content_268 = 64'h000000000000010c;
  assign content_269 = 64'h000000000000010d;
  assign content_270 = 64'h000000000000010e;
  assign content_271 = 64'h000000000000010f;
  assign content_272 = 64'h0000000000000110;
  assign content_273 = 64'h0000000000000111;
  assign content_274 = 64'h0000000000000112;
  assign content_275 = 64'h0000000000000113;
  assign content_276 = 64'h0000000000000114;
  assign content_277 = 64'h0000000000000115;
  assign content_278 = 64'h0000000000000116;
  assign content_279 = 64'h0000000000000117;
  assign content_280 = 64'h0000000000000118;
  assign content_281 = 64'h0000000000000119;
  assign content_282 = 64'h000000000000011a;
  assign content_283 = 64'h000000000000011b;
  assign content_284 = 64'h000000000000011c;
  assign content_285 = 64'h000000000000011d;
  assign content_286 = 64'h000000000000011e;
  assign content_287 = 64'h000000000000011f;
  assign content_288 = 64'h0000000000000120;
  assign content_289 = 64'h0000000000000121;
  assign content_290 = 64'h0000000000000122;
  assign content_291 = 64'h0000000000000123;
  assign content_292 = 64'h0000000000000124;
  assign content_293 = 64'h0000000000000125;
  assign content_294 = 64'h0000000000000126;
  assign content_295 = 64'h0000000000000127;
  assign content_296 = 64'h0000000000000128;
  assign content_297 = 64'h0000000000000129;
  assign content_298 = 64'h000000000000012a;
  assign content_299 = 64'h000000000000012b;
  assign content_300 = 64'h000000000000012c;
  assign content_301 = 64'h000000000000012d;
  assign content_302 = 64'h000000000000012e;
  assign content_303 = 64'h000000000000012f;
  assign content_304 = 64'h0000000000000130;
  assign content_305 = 64'h0000000000000131;
  assign content_306 = 64'h0000000000000132;
  assign content_307 = 64'h0000000000000133;
  assign content_308 = 64'h0000000000000134;
  assign content_309 = 64'h0000000000000135;
  assign content_310 = 64'h0000000000000136;
  assign content_311 = 64'h0000000000000137;
  assign content_312 = 64'h0000000000000138;
  assign content_313 = 64'h0000000000000139;
  assign content_314 = 64'h000000000000013a;
  assign content_315 = 64'h000000000000013b;
  assign content_316 = 64'h000000000000013c;
  assign content_317 = 64'h000000000000013d;
  assign content_318 = 64'h000000000000013e;
  assign content_319 = 64'h000000000000013f;
  assign content_320 = 64'h0000000000000140;
  assign content_321 = 64'h0000000000000141;
  assign content_322 = 64'h0000000000000142;
  assign content_323 = 64'h0000000000000143;
  assign content_324 = 64'h0000000000000144;
  assign content_325 = 64'h0000000000000145;
  assign content_326 = 64'h0000000000000146;
  assign content_327 = 64'h0000000000000147;
  assign content_328 = 64'h0000000000000148;
  assign content_329 = 64'h0000000000000149;
  assign content_330 = 64'h000000000000014a;
  assign content_331 = 64'h000000000000014b;
  assign content_332 = 64'h000000000000014c;
  assign content_333 = 64'h000000000000014d;
  assign content_334 = 64'h000000000000014e;
  assign content_335 = 64'h000000000000014f;
  assign content_336 = 64'h0000000000000150;
  assign content_337 = 64'h0000000000000151;
  assign content_338 = 64'h0000000000000152;
  assign content_339 = 64'h0000000000000153;
  assign content_340 = 64'h0000000000000154;
  assign content_341 = 64'h0000000000000155;
  assign content_342 = 64'h0000000000000156;
  assign content_343 = 64'h0000000000000157;
  assign content_344 = 64'h0000000000000158;
  assign content_345 = 64'h0000000000000159;
  assign content_346 = 64'h000000000000015a;
  assign content_347 = 64'h000000000000015b;
  assign content_348 = 64'h000000000000015c;
  assign content_349 = 64'h000000000000015d;
  assign content_350 = 64'h000000000000015e;
  assign content_351 = 64'h000000000000015f;
  assign content_352 = 64'h0000000000000160;
  assign content_353 = 64'h0000000000000161;
  assign content_354 = 64'h0000000000000162;
  assign content_355 = 64'h0000000000000163;
  assign content_356 = 64'h0000000000000164;
  assign content_357 = 64'h0000000000000165;
  assign content_358 = 64'h0000000000000166;
  assign content_359 = 64'h0000000000000167;
  assign content_360 = 64'h0000000000000168;
  assign content_361 = 64'h0000000000000169;
  assign content_362 = 64'h000000000000016a;
  assign content_363 = 64'h000000000000016b;
  assign content_364 = 64'h000000000000016c;
  assign content_365 = 64'h000000000000016d;
  assign content_366 = 64'h000000000000016e;
  assign content_367 = 64'h000000000000016f;
  assign content_368 = 64'h0000000000000170;
  assign content_369 = 64'h0000000000000171;
  assign content_370 = 64'h0000000000000172;
  assign content_371 = 64'h0000000000000173;
  assign content_372 = 64'h0000000000000174;
  assign content_373 = 64'h0000000000000175;
  assign content_374 = 64'h0000000000000176;
  assign content_375 = 64'h0000000000000177;
  assign content_376 = 64'h0000000000000178;
  assign content_377 = 64'h0000000000000179;
  assign content_378 = 64'h000000000000017a;
  assign content_379 = 64'h000000000000017b;
  assign content_380 = 64'h000000000000017c;
  assign content_381 = 64'h000000000000017d;
  assign content_382 = 64'h000000000000017e;
  assign content_383 = 64'h000000000000017f;
  assign content_384 = 64'h0000000000000180;
  assign content_385 = 64'h0000000000000181;
  assign content_386 = 64'h0000000000000182;
  assign content_387 = 64'h0000000000000183;
  assign content_388 = 64'h0000000000000184;
  assign content_389 = 64'h0000000000000185;
  assign content_390 = 64'h0000000000000186;
  assign content_391 = 64'h0000000000000187;
  assign content_392 = 64'h0000000000000188;
  assign content_393 = 64'h0000000000000189;
  assign content_394 = 64'h000000000000018a;
  assign content_395 = 64'h000000000000018b;
  assign content_396 = 64'h000000000000018c;
  assign content_397 = 64'h000000000000018d;
  assign content_398 = 64'h000000000000018e;
  assign content_399 = 64'h000000000000018f;
  assign content_400 = 64'h0000000000000190;
  assign content_401 = 64'h0000000000000191;
  assign content_402 = 64'h0000000000000192;
  assign content_403 = 64'h0000000000000193;
  assign content_404 = 64'h0000000000000194;
  assign content_405 = 64'h0000000000000195;
  assign content_406 = 64'h0000000000000196;
  assign content_407 = 64'h0000000000000197;
  assign content_408 = 64'h0000000000000198;
  assign content_409 = 64'h0000000000000199;
  assign content_410 = 64'h000000000000019a;
  assign content_411 = 64'h000000000000019b;
  assign content_412 = 64'h000000000000019c;
  assign content_413 = 64'h000000000000019d;
  assign content_414 = 64'h000000000000019e;
  assign content_415 = 64'h000000000000019f;
  assign content_416 = 64'h00000000000001a0;
  assign content_417 = 64'h00000000000001a1;
  assign content_418 = 64'h00000000000001a2;
  assign content_419 = 64'h00000000000001a3;
  assign content_420 = 64'h00000000000001a4;
  assign content_421 = 64'h00000000000001a5;
  assign content_422 = 64'h00000000000001a6;
  assign content_423 = 64'h00000000000001a7;
  assign content_424 = 64'h00000000000001a8;
  assign content_425 = 64'h00000000000001a9;
  assign content_426 = 64'h00000000000001aa;
  assign content_427 = 64'h00000000000001ab;
  assign content_428 = 64'h00000000000001ac;
  assign content_429 = 64'h00000000000001ad;
  assign content_430 = 64'h00000000000001ae;
  assign content_431 = 64'h00000000000001af;
  assign content_432 = 64'h00000000000001b0;
  assign content_433 = 64'h00000000000001b1;
  assign content_434 = 64'h00000000000001b2;
  assign content_435 = 64'h00000000000001b3;
  assign content_436 = 64'h00000000000001b4;
  assign content_437 = 64'h00000000000001b5;
  assign content_438 = 64'h00000000000001b6;
  assign content_439 = 64'h00000000000001b7;
  assign content_440 = 64'h00000000000001b8;
  assign content_441 = 64'h00000000000001b9;
  assign content_442 = 64'h00000000000001ba;
  assign content_443 = 64'h00000000000001bb;
  assign content_444 = 64'h00000000000001bc;
  assign content_445 = 64'h00000000000001bd;
  assign content_446 = 64'h00000000000001be;
  assign content_447 = 64'h00000000000001bf;
  assign content_448 = 64'h00000000000001c0;
  assign content_449 = 64'h00000000000001c1;
  assign content_450 = 64'h00000000000001c2;
  assign content_451 = 64'h00000000000001c3;
  assign content_452 = 64'h00000000000001c4;
  assign content_453 = 64'h00000000000001c5;
  assign content_454 = 64'h00000000000001c6;
  assign content_455 = 64'h00000000000001c7;
  assign content_456 = 64'h00000000000001c8;
  assign content_457 = 64'h00000000000001c9;
  assign content_458 = 64'h00000000000001ca;
  assign content_459 = 64'h00000000000001cb;
  assign content_460 = 64'h00000000000001cc;
  assign content_461 = 64'h00000000000001cd;
  assign content_462 = 64'h00000000000001ce;
  assign content_463 = 64'h00000000000001cf;
  assign content_464 = 64'h00000000000001d0;
  assign content_465 = 64'h00000000000001d1;
  assign content_466 = 64'h00000000000001d2;
  assign content_467 = 64'h00000000000001d3;
  assign content_468 = 64'h00000000000001d4;
  assign content_469 = 64'h00000000000001d5;
  assign content_470 = 64'h00000000000001d6;
  assign content_471 = 64'h00000000000001d7;
  assign content_472 = 64'h00000000000001d8;
  assign content_473 = 64'h00000000000001d9;
  assign content_474 = 64'h00000000000001da;
  assign content_475 = 64'h00000000000001db;
  assign content_476 = 64'h00000000000001dc;
  assign content_477 = 64'h00000000000001dd;
  assign content_478 = 64'h00000000000001de;
  assign content_479 = 64'h00000000000001df;
  assign content_480 = 64'h00000000000001e0;
  assign content_481 = 64'h00000000000001e1;
  assign content_482 = 64'h00000000000001e2;
  assign content_483 = 64'h00000000000001e3;
  assign content_484 = 64'h00000000000001e4;
  assign content_485 = 64'h00000000000001e5;
  assign content_486 = 64'h00000000000001e6;
  assign content_487 = 64'h00000000000001e7;
  assign content_488 = 64'h00000000000001e8;
  assign content_489 = 64'h00000000000001e9;
  assign content_490 = 64'h00000000000001ea;
  assign content_491 = 64'h00000000000001eb;
  assign content_492 = 64'h00000000000001ec;
  assign content_493 = 64'h00000000000001ed;
  assign content_494 = 64'h00000000000001ee;
  assign content_495 = 64'h00000000000001ef;
  assign content_496 = 64'h00000000000001f0;
  assign content_497 = 64'h00000000000001f1;
  assign content_498 = 64'h00000000000001f2;
  assign content_499 = 64'h00000000000001f3;
  assign content_500 = 64'h00000000000001f4;
  assign content_501 = 64'h00000000000001f5;
  assign content_502 = 64'h00000000000001f6;
  assign content_503 = 64'h00000000000001f7;
  assign content_504 = 64'h00000000000001f8;
  assign content_505 = 64'h00000000000001f9;
  assign content_506 = 64'h00000000000001fa;
  assign content_507 = 64'h00000000000001fb;
  assign content_508 = 64'h00000000000001fc;
  assign content_509 = 64'h00000000000001fd;
  assign content_510 = 64'h00000000000001fe;
  assign content_511 = 64'h00000000000001ff;
  assign content_512 = 64'h0000000000000200;
  assign content_513 = 64'h0000000000000201;
  assign content_514 = 64'h0000000000000202;
  assign content_515 = 64'h0000000000000203;
  assign content_516 = 64'h0000000000000204;
  assign content_517 = 64'h0000000000000205;
  assign content_518 = 64'h0000000000000206;
  assign content_519 = 64'h0000000000000207;
  assign content_520 = 64'h0000000000000208;
  assign content_521 = 64'h0000000000000209;
  assign content_522 = 64'h000000000000020a;
  assign content_523 = 64'h000000000000020b;
  assign content_524 = 64'h000000000000020c;
  assign content_525 = 64'h000000000000020d;
  assign content_526 = 64'h000000000000020e;
  assign content_527 = 64'h000000000000020f;
  assign content_528 = 64'h0000000000000210;
  assign content_529 = 64'h0000000000000211;
  assign content_530 = 64'h0000000000000212;
  assign content_531 = 64'h0000000000000213;
  assign content_532 = 64'h0000000000000214;
  assign content_533 = 64'h0000000000000215;
  assign content_534 = 64'h0000000000000216;
  assign content_535 = 64'h0000000000000217;
  assign content_536 = 64'h0000000000000218;
  assign content_537 = 64'h0000000000000219;
  assign content_538 = 64'h000000000000021a;
  assign content_539 = 64'h000000000000021b;
  assign content_540 = 64'h000000000000021c;
  assign content_541 = 64'h000000000000021d;
  assign content_542 = 64'h000000000000021e;
  assign content_543 = 64'h000000000000021f;
  assign content_544 = 64'h0000000000000220;
  assign content_545 = 64'h0000000000000221;
  assign content_546 = 64'h0000000000000222;
  assign content_547 = 64'h0000000000000223;
  assign content_548 = 64'h0000000000000224;
  assign content_549 = 64'h0000000000000225;
  assign content_550 = 64'h0000000000000226;
  assign content_551 = 64'h0000000000000227;
  assign content_552 = 64'h0000000000000228;
  assign content_553 = 64'h0000000000000229;
  assign content_554 = 64'h000000000000022a;
  assign content_555 = 64'h000000000000022b;
  assign content_556 = 64'h000000000000022c;
  assign content_557 = 64'h000000000000022d;
  assign content_558 = 64'h000000000000022e;
  assign content_559 = 64'h000000000000022f;
  assign content_560 = 64'h0000000000000230;
  assign content_561 = 64'h0000000000000231;
  assign content_562 = 64'h0000000000000232;
  assign content_563 = 64'h0000000000000233;
  assign content_564 = 64'h0000000000000234;
  assign content_565 = 64'h0000000000000235;
  assign content_566 = 64'h0000000000000236;
  assign content_567 = 64'h0000000000000237;
  assign content_568 = 64'h0000000000000238;
  assign content_569 = 64'h0000000000000239;
  assign content_570 = 64'h000000000000023a;
  assign content_571 = 64'h000000000000023b;
  assign content_572 = 64'h000000000000023c;
  assign content_573 = 64'h000000000000023d;
  assign content_574 = 64'h000000000000023e;
  assign content_575 = 64'h000000000000023f;
  assign content_576 = 64'h0000000000000240;
  assign content_577 = 64'h0000000000000241;
  assign content_578 = 64'h0000000000000242;
  assign content_579 = 64'h0000000000000243;
  assign content_580 = 64'h0000000000000244;
  assign content_581 = 64'h0000000000000245;
  assign content_582 = 64'h0000000000000246;
  assign content_583 = 64'h0000000000000247;
  assign content_584 = 64'h0000000000000248;
  assign content_585 = 64'h0000000000000249;
  assign content_586 = 64'h000000000000024a;
  assign content_587 = 64'h000000000000024b;
  assign content_588 = 64'h000000000000024c;
  assign content_589 = 64'h000000000000024d;
  assign content_590 = 64'h000000000000024e;
  assign content_591 = 64'h000000000000024f;
  assign content_592 = 64'h0000000000000250;
  assign content_593 = 64'h0000000000000251;
  assign content_594 = 64'h0000000000000252;
  assign content_595 = 64'h0000000000000253;
  assign content_596 = 64'h0000000000000254;
  assign content_597 = 64'h0000000000000255;
  assign content_598 = 64'h0000000000000256;
  assign content_599 = 64'h0000000000000257;
  assign content_600 = 64'h0000000000000258;
  assign content_601 = 64'h0000000000000259;
  assign content_602 = 64'h000000000000025a;
  assign content_603 = 64'h000000000000025b;
  assign content_604 = 64'h000000000000025c;
  assign content_605 = 64'h000000000000025d;
  assign content_606 = 64'h000000000000025e;
  assign content_607 = 64'h000000000000025f;
  assign content_608 = 64'h0000000000000260;
  assign content_609 = 64'h0000000000000261;
  assign content_610 = 64'h0000000000000262;
  assign content_611 = 64'h0000000000000263;
  assign content_612 = 64'h0000000000000264;
  assign content_613 = 64'h0000000000000265;
  assign content_614 = 64'h0000000000000266;
  assign content_615 = 64'h0000000000000267;
  assign content_616 = 64'h0000000000000268;
  assign content_617 = 64'h0000000000000269;
  assign content_618 = 64'h000000000000026a;
  assign content_619 = 64'h000000000000026b;
  assign content_620 = 64'h000000000000026c;
  assign content_621 = 64'h000000000000026d;
  assign content_622 = 64'h000000000000026e;
  assign content_623 = 64'h000000000000026f;
  assign content_624 = 64'h0000000000000270;
  assign content_625 = 64'h0000000000000271;
  assign content_626 = 64'h0000000000000272;
  assign content_627 = 64'h0000000000000273;
  assign content_628 = 64'h0000000000000274;
  assign content_629 = 64'h0000000000000275;
  assign content_630 = 64'h0000000000000276;
  assign content_631 = 64'h0000000000000277;
  assign content_632 = 64'h0000000000000278;
  assign content_633 = 64'h0000000000000279;
  assign content_634 = 64'h000000000000027a;
  assign content_635 = 64'h000000000000027b;
  assign content_636 = 64'h000000000000027c;
  assign content_637 = 64'h000000000000027d;
  assign content_638 = 64'h000000000000027e;
  assign content_639 = 64'h000000000000027f;
  assign content_640 = 64'h0000000000000280;
  assign content_641 = 64'h0000000000000281;
  assign content_642 = 64'h0000000000000282;
  assign content_643 = 64'h0000000000000283;
  assign content_644 = 64'h0000000000000284;
  assign content_645 = 64'h0000000000000285;
  assign content_646 = 64'h0000000000000286;
  assign content_647 = 64'h0000000000000287;
  assign content_648 = 64'h0000000000000288;
  assign content_649 = 64'h0000000000000289;
  assign content_650 = 64'h000000000000028a;
  assign content_651 = 64'h000000000000028b;
  assign content_652 = 64'h000000000000028c;
  assign content_653 = 64'h000000000000028d;
  assign content_654 = 64'h000000000000028e;
  assign content_655 = 64'h000000000000028f;
  assign content_656 = 64'h0000000000000290;
  assign content_657 = 64'h0000000000000291;
  assign content_658 = 64'h0000000000000292;
  assign content_659 = 64'h0000000000000293;
  assign content_660 = 64'h0000000000000294;
  assign content_661 = 64'h0000000000000295;
  assign content_662 = 64'h0000000000000296;
  assign content_663 = 64'h0000000000000297;
  assign content_664 = 64'h0000000000000298;
  assign content_665 = 64'h0000000000000299;
  assign content_666 = 64'h000000000000029a;
  assign content_667 = 64'h000000000000029b;
  assign content_668 = 64'h000000000000029c;
  assign content_669 = 64'h000000000000029d;
  assign content_670 = 64'h000000000000029e;
  assign content_671 = 64'h000000000000029f;
  assign content_672 = 64'h00000000000002a0;
  assign content_673 = 64'h00000000000002a1;
  assign content_674 = 64'h00000000000002a2;
  assign content_675 = 64'h00000000000002a3;
  assign content_676 = 64'h00000000000002a4;
  assign content_677 = 64'h00000000000002a5;
  assign content_678 = 64'h00000000000002a6;
  assign content_679 = 64'h00000000000002a7;
  assign content_680 = 64'h00000000000002a8;
  assign content_681 = 64'h00000000000002a9;
  assign content_682 = 64'h00000000000002aa;
  assign content_683 = 64'h00000000000002ab;
  assign content_684 = 64'h00000000000002ac;
  assign content_685 = 64'h00000000000002ad;
  assign content_686 = 64'h00000000000002ae;
  assign content_687 = 64'h00000000000002af;
  assign content_688 = 64'h00000000000002b0;
  assign content_689 = 64'h00000000000002b1;
  assign content_690 = 64'h00000000000002b2;
  assign content_691 = 64'h00000000000002b3;
  assign content_692 = 64'h00000000000002b4;
  assign content_693 = 64'h00000000000002b5;
  assign content_694 = 64'h00000000000002b6;
  assign content_695 = 64'h00000000000002b7;
  assign content_696 = 64'h00000000000002b8;
  assign content_697 = 64'h00000000000002b9;
  assign content_698 = 64'h00000000000002ba;
  assign content_699 = 64'h00000000000002bb;
  assign content_700 = 64'h00000000000002bc;
  assign content_701 = 64'h00000000000002bd;
  assign content_702 = 64'h00000000000002be;
  assign content_703 = 64'h00000000000002bf;
  assign content_704 = 64'h00000000000002c0;
  assign content_705 = 64'h00000000000002c1;
  assign content_706 = 64'h00000000000002c2;
  assign content_707 = 64'h00000000000002c3;
  assign content_708 = 64'h00000000000002c4;
  assign content_709 = 64'h00000000000002c5;
  assign content_710 = 64'h00000000000002c6;
  assign content_711 = 64'h00000000000002c7;
  assign content_712 = 64'h00000000000002c8;
  assign content_713 = 64'h00000000000002c9;
  assign content_714 = 64'h00000000000002ca;
  assign content_715 = 64'h00000000000002cb;
  assign content_716 = 64'h00000000000002cc;
  assign content_717 = 64'h00000000000002cd;
  assign content_718 = 64'h00000000000002ce;
  assign content_719 = 64'h00000000000002cf;
  assign content_720 = 64'h00000000000002d0;
  assign content_721 = 64'h00000000000002d1;
  assign content_722 = 64'h00000000000002d2;
  assign content_723 = 64'h00000000000002d3;
  assign content_724 = 64'h00000000000002d4;
  assign content_725 = 64'h00000000000002d5;
  assign content_726 = 64'h00000000000002d6;
  assign content_727 = 64'h00000000000002d7;
  assign content_728 = 64'h00000000000002d8;
  assign content_729 = 64'h00000000000002d9;
  assign content_730 = 64'h00000000000002da;
  assign content_731 = 64'h00000000000002db;
  assign content_732 = 64'h00000000000002dc;
  assign content_733 = 64'h00000000000002dd;
  assign content_734 = 64'h00000000000002de;
  assign content_735 = 64'h00000000000002df;
  assign content_736 = 64'h00000000000002e0;
  assign content_737 = 64'h00000000000002e1;
  assign content_738 = 64'h00000000000002e2;
  assign content_739 = 64'h00000000000002e3;
  assign content_740 = 64'h00000000000002e4;
  assign content_741 = 64'h00000000000002e5;
  assign content_742 = 64'h00000000000002e6;
  assign content_743 = 64'h00000000000002e7;
  assign content_744 = 64'h00000000000002e8;
  assign content_745 = 64'h00000000000002e9;
  assign content_746 = 64'h00000000000002ea;
  assign content_747 = 64'h00000000000002eb;
  assign content_748 = 64'h00000000000002ec;
  assign content_749 = 64'h00000000000002ed;
  assign content_750 = 64'h00000000000002ee;
  assign content_751 = 64'h00000000000002ef;
  assign content_752 = 64'h00000000000002f0;
  assign content_753 = 64'h00000000000002f1;
  assign content_754 = 64'h00000000000002f2;
  assign content_755 = 64'h00000000000002f3;
  assign content_756 = 64'h00000000000002f4;
  assign content_757 = 64'h00000000000002f5;
  assign content_758 = 64'h00000000000002f6;
  assign content_759 = 64'h00000000000002f7;
  assign content_760 = 64'h00000000000002f8;
  assign content_761 = 64'h00000000000002f9;
  assign content_762 = 64'h00000000000002fa;
  assign content_763 = 64'h00000000000002fb;
  assign content_764 = 64'h00000000000002fc;
  assign content_765 = 64'h00000000000002fd;
  assign content_766 = 64'h00000000000002fe;
  assign content_767 = 64'h00000000000002ff;
  assign content_768 = 64'h0000000000000300;
  assign content_769 = 64'h0000000000000301;
  assign content_770 = 64'h0000000000000302;
  assign content_771 = 64'h0000000000000303;
  assign content_772 = 64'h0000000000000304;
  assign content_773 = 64'h0000000000000305;
  assign content_774 = 64'h0000000000000306;
  assign content_775 = 64'h0000000000000307;
  assign content_776 = 64'h0000000000000308;
  assign content_777 = 64'h0000000000000309;
  assign content_778 = 64'h000000000000030a;
  assign content_779 = 64'h000000000000030b;
  assign content_780 = 64'h000000000000030c;
  assign content_781 = 64'h000000000000030d;
  assign content_782 = 64'h000000000000030e;
  assign content_783 = 64'h000000000000030f;
  assign content_784 = 64'h0000000000000310;
  assign content_785 = 64'h0000000000000311;
  assign content_786 = 64'h0000000000000312;
  assign content_787 = 64'h0000000000000313;
  assign content_788 = 64'h0000000000000314;
  assign content_789 = 64'h0000000000000315;
  assign content_790 = 64'h0000000000000316;
  assign content_791 = 64'h0000000000000317;
  assign content_792 = 64'h0000000000000318;
  assign content_793 = 64'h0000000000000319;
  assign content_794 = 64'h000000000000031a;
  assign content_795 = 64'h000000000000031b;
  assign content_796 = 64'h000000000000031c;
  assign content_797 = 64'h000000000000031d;
  assign content_798 = 64'h000000000000031e;
  assign content_799 = 64'h000000000000031f;
  assign content_800 = 64'h0000000000000320;
  assign content_801 = 64'h0000000000000321;
  assign content_802 = 64'h0000000000000322;
  assign content_803 = 64'h0000000000000323;
  assign content_804 = 64'h0000000000000324;
  assign content_805 = 64'h0000000000000325;
  assign content_806 = 64'h0000000000000326;
  assign content_807 = 64'h0000000000000327;
  assign content_808 = 64'h0000000000000328;
  assign content_809 = 64'h0000000000000329;
  assign content_810 = 64'h000000000000032a;
  assign content_811 = 64'h000000000000032b;
  assign content_812 = 64'h000000000000032c;
  assign content_813 = 64'h000000000000032d;
  assign content_814 = 64'h000000000000032e;
  assign content_815 = 64'h000000000000032f;
  assign content_816 = 64'h0000000000000330;
  assign content_817 = 64'h0000000000000331;
  assign content_818 = 64'h0000000000000332;
  assign content_819 = 64'h0000000000000333;
  assign content_820 = 64'h0000000000000334;
  assign content_821 = 64'h0000000000000335;
  assign content_822 = 64'h0000000000000336;
  assign content_823 = 64'h0000000000000337;
  assign content_824 = 64'h0000000000000338;
  assign content_825 = 64'h0000000000000339;
  assign content_826 = 64'h000000000000033a;
  assign content_827 = 64'h000000000000033b;
  assign content_828 = 64'h000000000000033c;
  assign content_829 = 64'h000000000000033d;
  assign content_830 = 64'h000000000000033e;
  assign content_831 = 64'h000000000000033f;
  assign content_832 = 64'h0000000000000340;
  assign content_833 = 64'h0000000000000341;
  assign content_834 = 64'h0000000000000342;
  assign content_835 = 64'h0000000000000343;
  assign content_836 = 64'h0000000000000344;
  assign content_837 = 64'h0000000000000345;
  assign content_838 = 64'h0000000000000346;
  assign content_839 = 64'h0000000000000347;
  assign content_840 = 64'h0000000000000348;
  assign content_841 = 64'h0000000000000349;
  assign content_842 = 64'h000000000000034a;
  assign content_843 = 64'h000000000000034b;
  assign content_844 = 64'h000000000000034c;
  assign content_845 = 64'h000000000000034d;
  assign content_846 = 64'h000000000000034e;
  assign content_847 = 64'h000000000000034f;
  assign content_848 = 64'h0000000000000350;
  assign content_849 = 64'h0000000000000351;
  assign content_850 = 64'h0000000000000352;
  assign content_851 = 64'h0000000000000353;
  assign content_852 = 64'h0000000000000354;
  assign content_853 = 64'h0000000000000355;
  assign content_854 = 64'h0000000000000356;
  assign content_855 = 64'h0000000000000357;
  assign content_856 = 64'h0000000000000358;
  assign content_857 = 64'h0000000000000359;
  assign content_858 = 64'h000000000000035a;
  assign content_859 = 64'h000000000000035b;
  assign content_860 = 64'h000000000000035c;
  assign content_861 = 64'h000000000000035d;
  assign content_862 = 64'h000000000000035e;
  assign content_863 = 64'h000000000000035f;
  assign content_864 = 64'h0000000000000360;
  assign content_865 = 64'h0000000000000361;
  assign content_866 = 64'h0000000000000362;
  assign content_867 = 64'h0000000000000363;
  assign content_868 = 64'h0000000000000364;
  assign content_869 = 64'h0000000000000365;
  assign content_870 = 64'h0000000000000366;
  assign content_871 = 64'h0000000000000367;
  assign content_872 = 64'h0000000000000368;
  assign content_873 = 64'h0000000000000369;
  assign content_874 = 64'h000000000000036a;
  assign content_875 = 64'h000000000000036b;
  assign content_876 = 64'h000000000000036c;
  assign content_877 = 64'h000000000000036d;
  assign content_878 = 64'h000000000000036e;
  assign content_879 = 64'h000000000000036f;
  assign content_880 = 64'h0000000000000370;
  assign content_881 = 64'h0000000000000371;
  assign content_882 = 64'h0000000000000372;
  assign content_883 = 64'h0000000000000373;
  assign content_884 = 64'h0000000000000374;
  assign content_885 = 64'h0000000000000375;
  assign content_886 = 64'h0000000000000376;
  assign content_887 = 64'h0000000000000377;
  assign content_888 = 64'h0000000000000378;
  assign content_889 = 64'h0000000000000379;
  assign content_890 = 64'h000000000000037a;
  assign content_891 = 64'h000000000000037b;
  assign content_892 = 64'h000000000000037c;
  assign content_893 = 64'h000000000000037d;
  assign content_894 = 64'h000000000000037e;
  assign content_895 = 64'h000000000000037f;
  assign content_896 = 64'h0000000000000380;
  assign content_897 = 64'h0000000000000381;
  assign content_898 = 64'h0000000000000382;
  assign content_899 = 64'h0000000000000383;
  assign content_900 = 64'h0000000000000384;
  assign content_901 = 64'h0000000000000385;
  assign content_902 = 64'h0000000000000386;
  assign content_903 = 64'h0000000000000387;
  assign content_904 = 64'h0000000000000388;
  assign content_905 = 64'h0000000000000389;
  assign content_906 = 64'h000000000000038a;
  assign content_907 = 64'h000000000000038b;
  assign content_908 = 64'h000000000000038c;
  assign content_909 = 64'h000000000000038d;
  assign content_910 = 64'h000000000000038e;
  assign content_911 = 64'h000000000000038f;
  assign content_912 = 64'h0000000000000390;
  assign content_913 = 64'h0000000000000391;
  assign content_914 = 64'h0000000000000392;
  assign content_915 = 64'h0000000000000393;
  assign content_916 = 64'h0000000000000394;
  assign content_917 = 64'h0000000000000395;
  assign content_918 = 64'h0000000000000396;
  assign content_919 = 64'h0000000000000397;
  assign content_920 = 64'h0000000000000398;
  assign content_921 = 64'h0000000000000399;
  assign content_922 = 64'h000000000000039a;
  assign content_923 = 64'h000000000000039b;
  assign content_924 = 64'h000000000000039c;
  assign content_925 = 64'h000000000000039d;
  assign content_926 = 64'h000000000000039e;
  assign content_927 = 64'h000000000000039f;
  assign content_928 = 64'h00000000000003a0;
  assign content_929 = 64'h00000000000003a1;
  assign content_930 = 64'h00000000000003a2;
  assign content_931 = 64'h00000000000003a3;
  assign content_932 = 64'h00000000000003a4;
  assign content_933 = 64'h00000000000003a5;
  assign content_934 = 64'h00000000000003a6;
  assign content_935 = 64'h00000000000003a7;
  assign content_936 = 64'h00000000000003a8;
  assign content_937 = 64'h00000000000003a9;
  assign content_938 = 64'h00000000000003aa;
  assign content_939 = 64'h00000000000003ab;
  assign content_940 = 64'h00000000000003ac;
  assign content_941 = 64'h00000000000003ad;
  assign content_942 = 64'h00000000000003ae;
  assign content_943 = 64'h00000000000003af;
  assign content_944 = 64'h00000000000003b0;
  assign content_945 = 64'h00000000000003b1;
  assign content_946 = 64'h00000000000003b2;
  assign content_947 = 64'h00000000000003b3;
  assign content_948 = 64'h00000000000003b4;
  assign content_949 = 64'h00000000000003b5;
  assign content_950 = 64'h00000000000003b6;
  assign content_951 = 64'h00000000000003b7;
  assign content_952 = 64'h00000000000003b8;
  assign content_953 = 64'h00000000000003b9;
  assign content_954 = 64'h00000000000003ba;
  assign content_955 = 64'h00000000000003bb;
  assign content_956 = 64'h00000000000003bc;
  assign content_957 = 64'h00000000000003bd;
  assign content_958 = 64'h00000000000003be;
  assign content_959 = 64'h00000000000003bf;
  assign content_960 = 64'h00000000000003c0;
  assign content_961 = 64'h00000000000003c1;
  assign content_962 = 64'h00000000000003c2;
  assign content_963 = 64'h00000000000003c3;
  assign content_964 = 64'h00000000000003c4;
  assign content_965 = 64'h00000000000003c5;
  assign content_966 = 64'h00000000000003c6;
  assign content_967 = 64'h00000000000003c7;
  assign content_968 = 64'h00000000000003c8;
  assign content_969 = 64'h00000000000003c9;
  assign content_970 = 64'h00000000000003ca;
  assign content_971 = 64'h00000000000003cb;
  assign content_972 = 64'h00000000000003cc;
  assign content_973 = 64'h00000000000003cd;
  assign content_974 = 64'h00000000000003ce;
  assign content_975 = 64'h00000000000003cf;
  assign content_976 = 64'h00000000000003d0;
  assign content_977 = 64'h00000000000003d1;
  assign content_978 = 64'h00000000000003d2;
  assign content_979 = 64'h00000000000003d3;
  assign content_980 = 64'h00000000000003d4;
  assign content_981 = 64'h00000000000003d5;
  assign content_982 = 64'h00000000000003d6;
  assign content_983 = 64'h00000000000003d7;
  assign content_984 = 64'h00000000000003d8;
  assign content_985 = 64'h00000000000003d9;
  assign content_986 = 64'h00000000000003da;
  assign content_987 = 64'h00000000000003db;
  assign content_988 = 64'h00000000000003dc;
  assign content_989 = 64'h00000000000003dd;
  assign content_990 = 64'h00000000000003de;
  assign content_991 = 64'h00000000000003df;
  assign content_992 = 64'h00000000000003e0;
  assign content_993 = 64'h00000000000003e1;
  assign content_994 = 64'h00000000000003e2;
  assign content_995 = 64'h00000000000003e3;
  assign content_996 = 64'h00000000000003e4;
  assign content_997 = 64'h00000000000003e5;
  assign content_998 = 64'h00000000000003e6;
  assign content_999 = 64'h00000000000003e7;
  assign content_1000 = 64'h00000000000003e8;
  assign content_1001 = 64'h00000000000003e9;
  assign content_1002 = 64'h00000000000003ea;
  assign content_1003 = 64'h00000000000003eb;
  assign content_1004 = 64'h00000000000003ec;
  assign content_1005 = 64'h00000000000003ed;
  assign content_1006 = 64'h00000000000003ee;
  assign content_1007 = 64'h00000000000003ef;
  assign content_1008 = 64'h00000000000003f0;
  assign content_1009 = 64'h00000000000003f1;
  assign content_1010 = 64'h00000000000003f2;
  assign content_1011 = 64'h00000000000003f3;
  assign content_1012 = 64'h00000000000003f4;
  assign content_1013 = 64'h00000000000003f5;
  assign content_1014 = 64'h00000000000003f6;
  assign content_1015 = 64'h00000000000003f7;
  assign content_1016 = 64'h00000000000003f8;
  assign content_1017 = 64'h00000000000003f9;
  assign content_1018 = 64'h00000000000003fa;
  assign content_1019 = 64'h00000000000003fb;
  assign content_1020 = 64'h00000000000003fc;
  assign content_1021 = 64'h00000000000003fd;
  assign content_1022 = 64'h00000000000003fe;
  assign content_1023 = 64'h00000000000003ff;
  assign _zz_1_ = (address >>> 3);
  always @ (*) begin
    if(memRead)begin
      readData = _zz_2_;
    end else begin
      readData = 64'h0;
    end
  end


endmodule
