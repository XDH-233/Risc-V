// Generator : SpinalHDL v1.4.0    git head : ecb5a80b713566f417ea3ea061f9969e73770a7f
// Date      : 17/07/2021, 08:18:14
// Component : instMem



module instMem (
  input      [8:0]    address,
  output     [31:0]   instruction 
);
  wire       [31:0]   _zz_2_;
  wire       [31:0]   inst_0;
  wire       [31:0]   inst_1;
  wire       [31:0]   inst_2;
  wire       [31:0]   inst_3;
  wire       [31:0]   inst_4;
  wire       [31:0]   inst_5;
  wire       [31:0]   inst_6;
  wire       [31:0]   inst_7;
  wire       [31:0]   inst_8;
  wire       [31:0]   inst_9;
  wire       [31:0]   inst_10;
  wire       [31:0]   inst_11;
  wire       [31:0]   inst_12;
  wire       [31:0]   inst_13;
  wire       [31:0]   inst_14;
  wire       [31:0]   inst_15;
  wire       [31:0]   inst_16;
  wire       [31:0]   inst_17;
  wire       [31:0]   inst_18;
  wire       [31:0]   inst_19;
  wire       [31:0]   inst_20;
  wire       [31:0]   inst_21;
  wire       [31:0]   inst_22;
  wire       [31:0]   inst_23;
  wire       [31:0]   inst_24;
  wire       [31:0]   inst_25;
  wire       [31:0]   inst_26;
  wire       [31:0]   inst_27;
  wire       [31:0]   inst_28;
  wire       [31:0]   inst_29;
  wire       [31:0]   inst_30;
  wire       [31:0]   inst_31;
  wire       [31:0]   inst_32;
  wire       [31:0]   inst_33;
  wire       [31:0]   inst_34;
  wire       [31:0]   inst_35;
  wire       [31:0]   inst_36;
  wire       [31:0]   inst_37;
  wire       [31:0]   inst_38;
  wire       [31:0]   inst_39;
  wire       [31:0]   inst_40;
  wire       [31:0]   inst_41;
  wire       [31:0]   inst_42;
  wire       [31:0]   inst_43;
  wire       [31:0]   inst_44;
  wire       [31:0]   inst_45;
  wire       [31:0]   inst_46;
  wire       [31:0]   inst_47;
  wire       [31:0]   inst_48;
  wire       [31:0]   inst_49;
  wire       [31:0]   inst_50;
  wire       [31:0]   inst_51;
  wire       [31:0]   inst_52;
  wire       [31:0]   inst_53;
  wire       [31:0]   inst_54;
  wire       [31:0]   inst_55;
  wire       [31:0]   inst_56;
  wire       [31:0]   inst_57;
  wire       [31:0]   inst_58;
  wire       [31:0]   inst_59;
  wire       [31:0]   inst_60;
  wire       [31:0]   inst_61;
  wire       [31:0]   inst_62;
  wire       [31:0]   inst_63;
  wire       [31:0]   inst_64;
  wire       [31:0]   inst_65;
  wire       [31:0]   inst_66;
  wire       [31:0]   inst_67;
  wire       [31:0]   inst_68;
  wire       [31:0]   inst_69;
  wire       [31:0]   inst_70;
  wire       [31:0]   inst_71;
  wire       [31:0]   inst_72;
  wire       [31:0]   inst_73;
  wire       [31:0]   inst_74;
  wire       [31:0]   inst_75;
  wire       [31:0]   inst_76;
  wire       [31:0]   inst_77;
  wire       [31:0]   inst_78;
  wire       [31:0]   inst_79;
  wire       [31:0]   inst_80;
  wire       [31:0]   inst_81;
  wire       [31:0]   inst_82;
  wire       [31:0]   inst_83;
  wire       [31:0]   inst_84;
  wire       [31:0]   inst_85;
  wire       [31:0]   inst_86;
  wire       [31:0]   inst_87;
  wire       [31:0]   inst_88;
  wire       [31:0]   inst_89;
  wire       [31:0]   inst_90;
  wire       [31:0]   inst_91;
  wire       [31:0]   inst_92;
  wire       [31:0]   inst_93;
  wire       [31:0]   inst_94;
  wire       [31:0]   inst_95;
  wire       [31:0]   inst_96;
  wire       [31:0]   inst_97;
  wire       [31:0]   inst_98;
  wire       [31:0]   inst_99;
  wire       [31:0]   inst_100;
  wire       [31:0]   inst_101;
  wire       [31:0]   inst_102;
  wire       [31:0]   inst_103;
  wire       [31:0]   inst_104;
  wire       [31:0]   inst_105;
  wire       [31:0]   inst_106;
  wire       [31:0]   inst_107;
  wire       [31:0]   inst_108;
  wire       [31:0]   inst_109;
  wire       [31:0]   inst_110;
  wire       [31:0]   inst_111;
  wire       [31:0]   inst_112;
  wire       [31:0]   inst_113;
  wire       [31:0]   inst_114;
  wire       [31:0]   inst_115;
  wire       [31:0]   inst_116;
  wire       [31:0]   inst_117;
  wire       [31:0]   inst_118;
  wire       [31:0]   inst_119;
  wire       [31:0]   inst_120;
  wire       [31:0]   inst_121;
  wire       [31:0]   inst_122;
  wire       [31:0]   inst_123;
  wire       [31:0]   inst_124;
  wire       [31:0]   inst_125;
  wire       [31:0]   inst_126;
  wire       [31:0]   inst_127;
  wire       [6:0]    _zz_1_;
  reg [31:0] mem [0:127];

  initial begin
    $readmemb("instMem.v_toplevel_mem.bin",mem);
  end
  assign _zz_2_ = mem[_zz_1_];
  assign inst_0 = 32'h0;
  assign inst_1 = 32'h0;
  assign inst_2 = 32'h00003083;
  assign inst_3 = 32'h00803103;
  assign inst_4 = 32'h01003183;
  assign inst_5 = 32'h00310233;
  assign inst_6 = 32'h0;
  assign inst_7 = 32'h0;
  assign inst_8 = 32'h0;
  assign inst_9 = 32'h0;
  assign inst_10 = 32'h0;
  assign inst_11 = 32'h0;
  assign inst_12 = 32'h0;
  assign inst_13 = 32'h0;
  assign inst_14 = 32'h0;
  assign inst_15 = 32'h0;
  assign inst_16 = 32'h0;
  assign inst_17 = 32'h0;
  assign inst_18 = 32'h0;
  assign inst_19 = 32'h0;
  assign inst_20 = 32'h0;
  assign inst_21 = 32'h0;
  assign inst_22 = 32'h0;
  assign inst_23 = 32'h0;
  assign inst_24 = 32'h0;
  assign inst_25 = 32'h0;
  assign inst_26 = 32'h0;
  assign inst_27 = 32'h0;
  assign inst_28 = 32'h0;
  assign inst_29 = 32'h0;
  assign inst_30 = 32'h0;
  assign inst_31 = 32'h0;
  assign inst_32 = 32'h0;
  assign inst_33 = 32'h0;
  assign inst_34 = 32'h0;
  assign inst_35 = 32'h0;
  assign inst_36 = 32'h0;
  assign inst_37 = 32'h0;
  assign inst_38 = 32'h0;
  assign inst_39 = 32'h0;
  assign inst_40 = 32'h0;
  assign inst_41 = 32'h0;
  assign inst_42 = 32'h0;
  assign inst_43 = 32'h0;
  assign inst_44 = 32'h0;
  assign inst_45 = 32'h0;
  assign inst_46 = 32'h0;
  assign inst_47 = 32'h0;
  assign inst_48 = 32'h0;
  assign inst_49 = 32'h0;
  assign inst_50 = 32'h0;
  assign inst_51 = 32'h0;
  assign inst_52 = 32'h0;
  assign inst_53 = 32'h0;
  assign inst_54 = 32'h0;
  assign inst_55 = 32'h0;
  assign inst_56 = 32'h0;
  assign inst_57 = 32'h0;
  assign inst_58 = 32'h0;
  assign inst_59 = 32'h0;
  assign inst_60 = 32'h0;
  assign inst_61 = 32'h0;
  assign inst_62 = 32'h0;
  assign inst_63 = 32'h0;
  assign inst_64 = 32'h0;
  assign inst_65 = 32'h0;
  assign inst_66 = 32'h0;
  assign inst_67 = 32'h0;
  assign inst_68 = 32'h0;
  assign inst_69 = 32'h0;
  assign inst_70 = 32'h0;
  assign inst_71 = 32'h0;
  assign inst_72 = 32'h0;
  assign inst_73 = 32'h0;
  assign inst_74 = 32'h0;
  assign inst_75 = 32'h0;
  assign inst_76 = 32'h0;
  assign inst_77 = 32'h0;
  assign inst_78 = 32'h0;
  assign inst_79 = 32'h0;
  assign inst_80 = 32'h0;
  assign inst_81 = 32'h0;
  assign inst_82 = 32'h0;
  assign inst_83 = 32'h0;
  assign inst_84 = 32'h0;
  assign inst_85 = 32'h0;
  assign inst_86 = 32'h0;
  assign inst_87 = 32'h0;
  assign inst_88 = 32'h0;
  assign inst_89 = 32'h0;
  assign inst_90 = 32'h0;
  assign inst_91 = 32'h0;
  assign inst_92 = 32'h0;
  assign inst_93 = 32'h0;
  assign inst_94 = 32'h0;
  assign inst_95 = 32'h0;
  assign inst_96 = 32'h0;
  assign inst_97 = 32'h0;
  assign inst_98 = 32'h0;
  assign inst_99 = 32'h0;
  assign inst_100 = 32'h0;
  assign inst_101 = 32'h0;
  assign inst_102 = 32'h0;
  assign inst_103 = 32'h0;
  assign inst_104 = 32'h0;
  assign inst_105 = 32'h0;
  assign inst_106 = 32'h0;
  assign inst_107 = 32'h0;
  assign inst_108 = 32'h0;
  assign inst_109 = 32'h0;
  assign inst_110 = 32'h0;
  assign inst_111 = 32'h0;
  assign inst_112 = 32'h0;
  assign inst_113 = 32'h0;
  assign inst_114 = 32'h0;
  assign inst_115 = 32'h0;
  assign inst_116 = 32'h0;
  assign inst_117 = 32'h0;
  assign inst_118 = 32'h0;
  assign inst_119 = 32'h0;
  assign inst_120 = 32'h0;
  assign inst_121 = 32'h0;
  assign inst_122 = 32'h0;
  assign inst_123 = 32'h0;
  assign inst_124 = 32'h0;
  assign inst_125 = 32'h0;
  assign inst_126 = 32'h0;
  assign inst_127 = 32'h0;
  assign _zz_1_ = (address >>> 2);
  assign instruction = _zz_2_;

endmodule
