// Generator : SpinalHDL v1.4.0    git head : ecb5a80b713566f417ea3ea061f9969e73770a7f
// Date      : 15/07/2021, 09:13:45
// Component : instMem



module instMem (
  input      [8:0]    address,
  output     [31:0]   instruction 
);
  wire       [31:0]   _zz_2_;
  wire       [31:0]   content_0;
  wire       [31:0]   content_1;
  wire       [31:0]   content_2;
  wire       [31:0]   content_3;
  wire       [31:0]   content_4;
  wire       [31:0]   content_5;
  wire       [31:0]   content_6;
  wire       [31:0]   content_7;
  wire       [31:0]   content_8;
  wire       [31:0]   content_9;
  wire       [31:0]   content_10;
  wire       [31:0]   content_11;
  wire       [31:0]   content_12;
  wire       [31:0]   content_13;
  wire       [31:0]   content_14;
  wire       [31:0]   content_15;
  wire       [31:0]   content_16;
  wire       [31:0]   content_17;
  wire       [31:0]   content_18;
  wire       [31:0]   content_19;
  wire       [31:0]   content_20;
  wire       [31:0]   content_21;
  wire       [31:0]   content_22;
  wire       [31:0]   content_23;
  wire       [31:0]   content_24;
  wire       [31:0]   content_25;
  wire       [31:0]   content_26;
  wire       [31:0]   content_27;
  wire       [31:0]   content_28;
  wire       [31:0]   content_29;
  wire       [31:0]   content_30;
  wire       [31:0]   content_31;
  wire       [31:0]   content_32;
  wire       [31:0]   content_33;
  wire       [31:0]   content_34;
  wire       [31:0]   content_35;
  wire       [31:0]   content_36;
  wire       [31:0]   content_37;
  wire       [31:0]   content_38;
  wire       [31:0]   content_39;
  wire       [31:0]   content_40;
  wire       [31:0]   content_41;
  wire       [31:0]   content_42;
  wire       [31:0]   content_43;
  wire       [31:0]   content_44;
  wire       [31:0]   content_45;
  wire       [31:0]   content_46;
  wire       [31:0]   content_47;
  wire       [31:0]   content_48;
  wire       [31:0]   content_49;
  wire       [31:0]   content_50;
  wire       [31:0]   content_51;
  wire       [31:0]   content_52;
  wire       [31:0]   content_53;
  wire       [31:0]   content_54;
  wire       [31:0]   content_55;
  wire       [31:0]   content_56;
  wire       [31:0]   content_57;
  wire       [31:0]   content_58;
  wire       [31:0]   content_59;
  wire       [31:0]   content_60;
  wire       [31:0]   content_61;
  wire       [31:0]   content_62;
  wire       [31:0]   content_63;
  wire       [31:0]   content_64;
  wire       [31:0]   content_65;
  wire       [31:0]   content_66;
  wire       [31:0]   content_67;
  wire       [31:0]   content_68;
  wire       [31:0]   content_69;
  wire       [31:0]   content_70;
  wire       [31:0]   content_71;
  wire       [31:0]   content_72;
  wire       [31:0]   content_73;
  wire       [31:0]   content_74;
  wire       [31:0]   content_75;
  wire       [31:0]   content_76;
  wire       [31:0]   content_77;
  wire       [31:0]   content_78;
  wire       [31:0]   content_79;
  wire       [31:0]   content_80;
  wire       [31:0]   content_81;
  wire       [31:0]   content_82;
  wire       [31:0]   content_83;
  wire       [31:0]   content_84;
  wire       [31:0]   content_85;
  wire       [31:0]   content_86;
  wire       [31:0]   content_87;
  wire       [31:0]   content_88;
  wire       [31:0]   content_89;
  wire       [31:0]   content_90;
  wire       [31:0]   content_91;
  wire       [31:0]   content_92;
  wire       [31:0]   content_93;
  wire       [31:0]   content_94;
  wire       [31:0]   content_95;
  wire       [31:0]   content_96;
  wire       [31:0]   content_97;
  wire       [31:0]   content_98;
  wire       [31:0]   content_99;
  wire       [31:0]   content_100;
  wire       [31:0]   content_101;
  wire       [31:0]   content_102;
  wire       [31:0]   content_103;
  wire       [31:0]   content_104;
  wire       [31:0]   content_105;
  wire       [31:0]   content_106;
  wire       [31:0]   content_107;
  wire       [31:0]   content_108;
  wire       [31:0]   content_109;
  wire       [31:0]   content_110;
  wire       [31:0]   content_111;
  wire       [31:0]   content_112;
  wire       [31:0]   content_113;
  wire       [31:0]   content_114;
  wire       [31:0]   content_115;
  wire       [31:0]   content_116;
  wire       [31:0]   content_117;
  wire       [31:0]   content_118;
  wire       [31:0]   content_119;
  wire       [31:0]   content_120;
  wire       [31:0]   content_121;
  wire       [31:0]   content_122;
  wire       [31:0]   content_123;
  wire       [31:0]   content_124;
  wire       [31:0]   content_125;
  wire       [31:0]   content_126;
  wire       [31:0]   content_127;
  wire       [6:0]    _zz_1_;
  reg [31:0] mem [0:127];

  initial begin
    $readmemb("instMem.v_toplevel_mem.bin",mem);
  end
  assign _zz_2_ = mem[_zz_1_];
  assign content_0 = 32'h0;
  assign content_1 = 32'h00000001;
  assign content_2 = 32'h00000002;
  assign content_3 = 32'h00000003;
  assign content_4 = 32'h00000004;
  assign content_5 = 32'h00000005;
  assign content_6 = 32'h00000006;
  assign content_7 = 32'h00000007;
  assign content_8 = 32'h00000008;
  assign content_9 = 32'h00000009;
  assign content_10 = 32'h0000000a;
  assign content_11 = 32'h0000000b;
  assign content_12 = 32'h0000000c;
  assign content_13 = 32'h0000000d;
  assign content_14 = 32'h0000000e;
  assign content_15 = 32'h0000000f;
  assign content_16 = 32'h00000010;
  assign content_17 = 32'h00000011;
  assign content_18 = 32'h00000012;
  assign content_19 = 32'h00000013;
  assign content_20 = 32'h00000014;
  assign content_21 = 32'h00000015;
  assign content_22 = 32'h00000016;
  assign content_23 = 32'h00000017;
  assign content_24 = 32'h00000018;
  assign content_25 = 32'h00000019;
  assign content_26 = 32'h0000001a;
  assign content_27 = 32'h0000001b;
  assign content_28 = 32'h0000001c;
  assign content_29 = 32'h0000001d;
  assign content_30 = 32'h0000001e;
  assign content_31 = 32'h0000001f;
  assign content_32 = 32'h00000020;
  assign content_33 = 32'h00000021;
  assign content_34 = 32'h00000022;
  assign content_35 = 32'h00000023;
  assign content_36 = 32'h00000024;
  assign content_37 = 32'h00000025;
  assign content_38 = 32'h00000026;
  assign content_39 = 32'h00000027;
  assign content_40 = 32'h00000028;
  assign content_41 = 32'h00000029;
  assign content_42 = 32'h0000002a;
  assign content_43 = 32'h0000002b;
  assign content_44 = 32'h0000002c;
  assign content_45 = 32'h0000002d;
  assign content_46 = 32'h0000002e;
  assign content_47 = 32'h0000002f;
  assign content_48 = 32'h00000030;
  assign content_49 = 32'h00000031;
  assign content_50 = 32'h00000032;
  assign content_51 = 32'h00000033;
  assign content_52 = 32'h00000034;
  assign content_53 = 32'h00000035;
  assign content_54 = 32'h00000036;
  assign content_55 = 32'h00000037;
  assign content_56 = 32'h00000038;
  assign content_57 = 32'h00000039;
  assign content_58 = 32'h0000003a;
  assign content_59 = 32'h0000003b;
  assign content_60 = 32'h0000003c;
  assign content_61 = 32'h0000003d;
  assign content_62 = 32'h0000003e;
  assign content_63 = 32'h0000003f;
  assign content_64 = 32'h00000040;
  assign content_65 = 32'h00000041;
  assign content_66 = 32'h00000042;
  assign content_67 = 32'h00000043;
  assign content_68 = 32'h00000044;
  assign content_69 = 32'h00000045;
  assign content_70 = 32'h00000046;
  assign content_71 = 32'h00000047;
  assign content_72 = 32'h00000048;
  assign content_73 = 32'h00000049;
  assign content_74 = 32'h0000004a;
  assign content_75 = 32'h0000004b;
  assign content_76 = 32'h0000004c;
  assign content_77 = 32'h0000004d;
  assign content_78 = 32'h0000004e;
  assign content_79 = 32'h0000004f;
  assign content_80 = 32'h00000050;
  assign content_81 = 32'h00000051;
  assign content_82 = 32'h00000052;
  assign content_83 = 32'h00000053;
  assign content_84 = 32'h00000054;
  assign content_85 = 32'h00000055;
  assign content_86 = 32'h00000056;
  assign content_87 = 32'h00000057;
  assign content_88 = 32'h00000058;
  assign content_89 = 32'h00000059;
  assign content_90 = 32'h0000005a;
  assign content_91 = 32'h0000005b;
  assign content_92 = 32'h0000005c;
  assign content_93 = 32'h0000005d;
  assign content_94 = 32'h0000005e;
  assign content_95 = 32'h0000005f;
  assign content_96 = 32'h00000060;
  assign content_97 = 32'h00000061;
  assign content_98 = 32'h00000062;
  assign content_99 = 32'h00000063;
  assign content_100 = 32'h00000064;
  assign content_101 = 32'h00000065;
  assign content_102 = 32'h00000066;
  assign content_103 = 32'h00000067;
  assign content_104 = 32'h00000068;
  assign content_105 = 32'h00000069;
  assign content_106 = 32'h0000006a;
  assign content_107 = 32'h0000006b;
  assign content_108 = 32'h0000006c;
  assign content_109 = 32'h0000006d;
  assign content_110 = 32'h0000006e;
  assign content_111 = 32'h0000006f;
  assign content_112 = 32'h00000070;
  assign content_113 = 32'h00000071;
  assign content_114 = 32'h00000072;
  assign content_115 = 32'h00000073;
  assign content_116 = 32'h00000074;
  assign content_117 = 32'h00000075;
  assign content_118 = 32'h00000076;
  assign content_119 = 32'h00000077;
  assign content_120 = 32'h00000078;
  assign content_121 = 32'h00000079;
  assign content_122 = 32'h0000007a;
  assign content_123 = 32'h0000007b;
  assign content_124 = 32'h0000007c;
  assign content_125 = 32'h0000007d;
  assign content_126 = 32'h0000007e;
  assign content_127 = 32'h0000007f;
  assign _zz_1_ = (address >>> 2);
  assign instruction = _zz_2_;

endmodule
